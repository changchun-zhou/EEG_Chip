# Created by MC2 : Version 2006.09.01.d on 2024/04/08, 13:49:31

###############################################################################
#        Software       : TSMC MEMORY COMPILER 2006.09.01.d
#        Technology     : 65 nm CMOS LOGIC Low Power LowK Cu 1P9M 1.2
#                         Mix-vt logic, High-vt SRAM
#        Memory Type    : TSMC 65nm low power SP SRAM Without Redundancy
#        Library Name   : ts1n65lpa1024x4m4
#        Library Version: 140a
#        Generated Time : 2024/04/08, 13:49:29
###############################################################################
#
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
#
###############################################################################
 
MACRO TS1N65LPA1024X4M4
	CLASS BLOCK ;
	FOREIGN TS1N65LPA1024X4M4 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 62.445 BY 181.555 ;
	SYMMETRY X Y R90 ;

	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 33.395 0.000 33.915 0.520 ;
			LAYER M3 ;
			RECT 33.395 0.000 33.915 0.520 ;
			LAYER M1 ;
			RECT 33.395 0.000 33.915 0.520 ;
		END
	END A[0]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 35.995 0.000 36.515 0.520 ;
			LAYER M3 ;
			RECT 35.995 0.000 36.515 0.520 ;
			LAYER M1 ;
			RECT 35.995 0.000 36.515 0.520 ;
		END
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 32.310 0.000 32.830 0.520 ;
			LAYER M1 ;
			RECT 32.310 0.000 32.830 0.520 ;
			LAYER M2 ;
			RECT 32.310 0.000 32.830 0.520 ;
		END
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 30.430 0.000 30.950 0.520 ;
			LAYER M2 ;
			RECT 30.430 0.000 30.950 0.520 ;
			LAYER M3 ;
			RECT 30.430 0.000 30.950 0.520 ;
		END
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 26.670 0.000 27.190 0.520 ;
			LAYER M1 ;
			RECT 26.670 0.000 27.190 0.520 ;
			LAYER M2 ;
			RECT 26.670 0.000 27.190 0.520 ;
		END
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 24.790 0.000 25.310 0.520 ;
			LAYER M1 ;
			RECT 24.790 0.000 25.310 0.520 ;
			LAYER M3 ;
			RECT 24.790 0.000 25.310 0.520 ;
		END
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 22.910 0.000 23.430 0.520 ;
			LAYER M2 ;
			RECT 22.910 0.000 23.430 0.520 ;
			LAYER M3 ;
			RECT 22.910 0.000 23.430 0.520 ;
		END
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 19.150 0.000 19.670 0.520 ;
			LAYER M3 ;
			RECT 19.150 0.000 19.670 0.520 ;
			LAYER M2 ;
			RECT 19.150 0.000 19.670 0.520 ;
		END
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 17.270 0.000 17.790 0.520 ;
			LAYER M1 ;
			RECT 17.270 0.000 17.790 0.520 ;
			LAYER M3 ;
			RECT 17.270 0.000 17.790 0.520 ;
		END
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 15.390 0.000 15.910 0.520 ;
			LAYER M2 ;
			RECT 15.390 0.000 15.910 0.520 ;
			LAYER M3 ;
			RECT 15.390 0.000 15.910 0.520 ;
		END
	END A[9]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 5.250 0.000 5.770 0.520 ;
			LAYER M1 ;
			RECT 5.250 0.000 5.770 0.520 ;
			LAYER M3 ;
			RECT 5.250 0.000 5.770 0.520 ;
		END
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 9.450 0.000 9.970 0.520 ;
			LAYER M3 ;
			RECT 9.450 0.000 9.970 0.520 ;
			LAYER M2 ;
			RECT 9.450 0.000 9.970 0.520 ;
		END
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 52.475 0.000 52.995 0.520 ;
			LAYER M1 ;
			RECT 52.475 0.000 52.995 0.520 ;
			LAYER M3 ;
			RECT 52.475 0.000 52.995 0.520 ;
		END
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 56.675 0.000 57.195 0.520 ;
			LAYER M1 ;
			RECT 56.675 0.000 57.195 0.520 ;
			LAYER M3 ;
			RECT 56.675 0.000 57.195 0.520 ;
		END
	END BWEB[3]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 41.240 0.000 41.760 0.520 ;
			LAYER M3 ;
			RECT 41.240 0.000 41.760 0.520 ;
			LAYER M2 ;
			RECT 41.240 0.000 41.760 0.520 ;
		END
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 47.670 0.000 48.190 0.520 ;
			LAYER M3 ;
			RECT 47.670 0.000 48.190 0.520 ;
			LAYER M1 ;
			RECT 47.670 0.000 48.190 0.520 ;
		END
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 1.970 0.000 2.490 0.520 ;
			LAYER M2 ;
			RECT 1.970 0.000 2.490 0.520 ;
			LAYER M3 ;
			RECT 1.970 0.000 2.490 0.520 ;
		END
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 6.170 0.000 6.690 0.520 ;
			LAYER M2 ;
			RECT 6.170 0.000 6.690 0.520 ;
			LAYER M1 ;
			RECT 6.170 0.000 6.690 0.520 ;
		END
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 55.755 0.000 56.275 0.520 ;
			LAYER M1 ;
			RECT 55.755 0.000 56.275 0.520 ;
			LAYER M2 ;
			RECT 55.755 0.000 56.275 0.520 ;
		END
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 59.955 0.000 60.475 0.520 ;
			LAYER M2 ;
			RECT 59.955 0.000 60.475 0.520 ;
			LAYER M3 ;
			RECT 59.955 0.000 60.475 0.520 ;
		END
	END D[3]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 3.610 0.000 4.130 0.520 ;
			LAYER M3 ;
			RECT 3.610 0.000 4.130 0.520 ;
			LAYER M1 ;
			RECT 3.610 0.000 4.130 0.520 ;
		END
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 7.810 0.000 8.330 0.520 ;
			LAYER M1 ;
			RECT 7.810 0.000 8.330 0.520 ;
			LAYER M3 ;
			RECT 7.810 0.000 8.330 0.520 ;
		END
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 54.115 0.000 54.635 0.520 ;
			LAYER M2 ;
			RECT 54.115 0.000 54.635 0.520 ;
			LAYER M3 ;
			RECT 54.115 0.000 54.635 0.520 ;
		END
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 58.315 0.000 58.835 0.520 ;
			LAYER M2 ;
			RECT 58.315 0.000 58.835 0.520 ;
			LAYER M3 ;
			RECT 58.315 0.000 58.835 0.520 ;
		END
	END Q[3]

	PIN TSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 51.445 0.000 51.965 0.520 ;
			LAYER M3 ;
			RECT 51.445 0.000 51.965 0.520 ;
			LAYER M2 ;
			RECT 51.445 0.000 51.965 0.520 ;
		END
	END TSEL[0]

	PIN TSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 50.725 0.000 51.245 0.520 ;
			LAYER M3 ;
			RECT 50.725 0.000 51.245 0.520 ;
			LAYER M1 ;
			RECT 50.725 0.000 51.245 0.520 ;
		END
	END TSEL[1]

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 39.775 0.000 40.295 0.520 ;
			LAYER M1 ;
			RECT 39.775 0.000 40.295 0.520 ;
			LAYER M3 ;
			RECT 39.775 0.000 40.295 0.520 ;
		END
	END WEB
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M5 ;
			RECT 0.000 10.000 29.970 14.000 ;
			LAYER M5 ;
			RECT 41.750 10.000 62.445 14.000 ;
			LAYER M5 ;
			RECT 0.000 26.000 29.970 30.000 ;
			LAYER M5 ;
			RECT 41.750 26.000 62.445 30.000 ;
			LAYER M5 ;
			RECT 0.000 42.000 29.970 46.000 ;
			LAYER M5 ;
			RECT 41.750 42.000 62.445 46.000 ;
			LAYER M5 ;
			RECT 0.000 58.000 29.970 62.000 ;
			LAYER M5 ;
			RECT 41.750 58.000 62.445 62.000 ;
			LAYER M5 ;
			RECT 0.000 74.000 29.970 78.000 ;
			LAYER M5 ;
			RECT 41.750 74.000 62.445 78.000 ;
			LAYER M5 ;
			RECT 0.000 90.000 29.970 94.000 ;
			LAYER M5 ;
			RECT 41.750 90.000 62.445 94.000 ;
			LAYER M5 ;
			RECT 0.000 106.000 29.970 110.000 ;
			LAYER M5 ;
			RECT 41.750 106.000 62.445 110.000 ;
			LAYER M5 ;
			RECT 0.000 122.000 29.970 126.000 ;
			LAYER M5 ;
			RECT 41.750 122.000 62.445 126.000 ;
			LAYER M5 ;
			RECT 0.000 138.000 29.970 142.000 ;
			LAYER M5 ;
			RECT 41.750 138.000 62.445 142.000 ;
			LAYER M5 ;
			RECT 0.000 154.000 29.970 158.000 ;
			LAYER M5 ;
			RECT 41.750 154.000 62.445 158.000 ;
			LAYER M5 ;
			RECT 0.000 170.000 29.970 174.000 ;
			LAYER M5 ;
			RECT 41.750 170.000 62.445 174.000 ;
		LAYER M4 ;
		RECT 0.140 0.730 0.470 181.555 ;
		LAYER M4 ;
		RECT 1.580 0.730 1.960 181.555 ;
		LAYER M4 ;
		RECT 3.680 0.730 4.060 181.555 ;
		LAYER M4 ;
		RECT 5.780 0.730 6.160 181.555 ;
		LAYER M4 ;
		RECT 7.880 0.730 8.260 181.555 ;
		LAYER M4 ;
		RECT 9.980 0.730 10.360 181.555 ;
		LAYER M4 ;
		RECT 22.810 0.730 25.810 181.555 ;
		LAYER M4 ;
		RECT 34.310 0.730 36.310 181.555 ;
		LAYER M4 ;
		RECT 41.750 0.730 43.750 181.555 ;
		LAYER M4 ;
		RECT 49.985 0.730 50.365 181.555 ;
		LAYER M4 ;
		RECT 52.085 0.730 52.465 181.555 ;
		LAYER M4 ;
		RECT 54.185 0.730 54.565 181.555 ;
		LAYER M4 ;
		RECT 56.285 0.730 56.665 181.555 ;
		LAYER M4 ;
		RECT 58.385 0.730 58.765 181.555 ;
		LAYER M4 ;
		RECT 60.485 0.730 60.865 181.555 ;
		LAYER M4 ;
		RECT 61.975 0.730 62.305 181.555 ;
		END
	END VDD

	PIN GND
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M5 ;
			RECT 0.000 2.000 29.970 6.000 ;
			LAYER M5 ;
			RECT 41.750 2.000 62.445 6.000 ;
			LAYER M5 ;
			RECT 0.000 18.000 29.970 22.000 ;
			LAYER M5 ;
			RECT 41.750 18.000 62.445 22.000 ;
			LAYER M5 ;
			RECT 0.000 34.000 29.970 38.000 ;
			LAYER M5 ;
			RECT 41.750 34.000 62.445 38.000 ;
			LAYER M5 ;
			RECT 0.000 50.000 29.970 54.000 ;
			LAYER M5 ;
			RECT 41.750 50.000 62.445 54.000 ;
			LAYER M5 ;
			RECT 0.000 66.000 29.970 70.000 ;
			LAYER M5 ;
			RECT 41.750 66.000 62.445 70.000 ;
			LAYER M5 ;
			RECT 0.000 82.000 29.970 86.000 ;
			LAYER M5 ;
			RECT 41.750 82.000 62.445 86.000 ;
			LAYER M5 ;
			RECT 0.000 98.000 29.970 102.000 ;
			LAYER M5 ;
			RECT 41.750 98.000 62.445 102.000 ;
			LAYER M5 ;
			RECT 0.000 114.000 29.970 118.000 ;
			LAYER M5 ;
			RECT 41.750 114.000 62.445 118.000 ;
			LAYER M5 ;
			RECT 0.000 130.000 29.970 134.000 ;
			LAYER M5 ;
			RECT 41.750 130.000 62.445 134.000 ;
			LAYER M5 ;
			RECT 0.000 146.000 29.970 150.000 ;
			LAYER M5 ;
			RECT 41.750 146.000 62.445 150.000 ;
			LAYER M5 ;
			RECT 0.000 162.000 29.970 166.000 ;
			LAYER M5 ;
			RECT 41.750 162.000 62.445 166.000 ;
		LAYER M4 ;
		RECT 1.035 0.730 1.415 181.555 ;
		LAYER M4 ;
		RECT 2.530 0.730 3.110 181.555 ;
		LAYER M4 ;
		RECT 4.630 0.730 5.210 181.555 ;
		LAYER M4 ;
		RECT 6.730 0.730 7.310 181.555 ;
		LAYER M4 ;
		RECT 8.830 0.730 9.410 181.555 ;
		LAYER M4 ;
		RECT 10.525 0.730 10.905 181.555 ;
		LAYER M4 ;
		RECT 21.910 0.730 22.310 181.555 ;
		LAYER M4 ;
		RECT 27.270 0.730 29.970 181.555 ;
		LAYER M4 ;
		RECT 45.675 0.730 48.875 181.555 ;
		LAYER M4 ;
		RECT 49.440 0.730 49.820 181.555 ;
		LAYER M4 ;
		RECT 50.935 0.730 51.515 181.555 ;
		LAYER M4 ;
		RECT 53.035 0.730 53.615 181.555 ;
		LAYER M4 ;
		RECT 55.135 0.730 55.715 181.555 ;
		LAYER M4 ;
		RECT 57.235 0.730 57.815 181.555 ;
		LAYER M4 ;
		RECT 59.335 0.730 59.915 181.555 ;
		LAYER M4 ;
		RECT 61.030 0.730 61.410 181.555 ;
		END
	END GND

	OBS
		# Pmesh blockages
		LAYER M5 ;
		RECT 2.000 10.000 27.970 12.000 ;
		LAYER M5 ;
		RECT 43.750 10.000 60.445 12.000 ;
		LAYER M5 ;
		RECT 2.000 26.000 27.970 28.000 ;
		LAYER M5 ;
		RECT 43.750 26.000 60.445 28.000 ;
		LAYER M5 ;
		RECT 2.000 42.000 27.970 44.000 ;
		LAYER M5 ;
		RECT 43.750 42.000 60.445 44.000 ;
		LAYER M5 ;
		RECT 2.000 58.000 27.970 60.000 ;
		LAYER M5 ;
		RECT 43.750 58.000 60.445 60.000 ;
		LAYER M5 ;
		RECT 2.000 74.000 27.970 76.000 ;
		LAYER M5 ;
		RECT 43.750 74.000 60.445 76.000 ;
		LAYER M5 ;
		RECT 2.000 90.000 27.970 92.000 ;
		LAYER M5 ;
		RECT 43.750 90.000 60.445 92.000 ;
		LAYER M5 ;
		RECT 2.000 106.000 27.970 108.000 ;
		LAYER M5 ;
		RECT 43.750 106.000 60.445 108.000 ;
		LAYER M5 ;
		RECT 2.000 122.000 27.970 124.000 ;
		LAYER M5 ;
		RECT 43.750 122.000 60.445 124.000 ;
		LAYER M5 ;
		RECT 2.000 138.000 27.970 140.000 ;
		LAYER M5 ;
		RECT 43.750 138.000 60.445 140.000 ;
		LAYER M5 ;
		RECT 2.000 154.000 27.970 156.000 ;
		LAYER M5 ;
		RECT 43.750 154.000 60.445 156.000 ;
		LAYER M5 ;
		RECT 2.000 170.000 27.970 172.000 ;
		LAYER M5 ;
		RECT 43.750 170.000 60.445 172.000 ;
		LAYER M5 ;
		RECT 2.000 2.000 27.970 4.000 ;
		LAYER M5 ;
		RECT 43.750 2.000 60.445 4.000 ;
		LAYER M5 ;
		RECT 2.000 18.000 27.970 20.000 ;
		LAYER M5 ;
		RECT 43.750 18.000 60.445 20.000 ;
		LAYER M5 ;
		RECT 2.000 34.000 27.970 36.000 ;
		LAYER M5 ;
		RECT 43.750 34.000 60.445 36.000 ;
		LAYER M5 ;
		RECT 2.000 50.000 27.970 52.000 ;
		LAYER M5 ;
		RECT 43.750 50.000 60.445 52.000 ;
		LAYER M5 ;
		RECT 2.000 66.000 27.970 68.000 ;
		LAYER M5 ;
		RECT 43.750 66.000 60.445 68.000 ;
		LAYER M5 ;
		RECT 2.000 82.000 27.970 84.000 ;
		LAYER M5 ;
		RECT 43.750 82.000 60.445 84.000 ;
		LAYER M5 ;
		RECT 2.000 98.000 27.970 100.000 ;
		LAYER M5 ;
		RECT 43.750 98.000 60.445 100.000 ;
		LAYER M5 ;
		RECT 2.000 114.000 27.970 116.000 ;
		LAYER M5 ;
		RECT 43.750 114.000 60.445 116.000 ;
		LAYER M5 ;
		RECT 2.000 130.000 27.970 132.000 ;
		LAYER M5 ;
		RECT 43.750 130.000 60.445 132.000 ;
		LAYER M5 ;
		RECT 2.000 146.000 27.970 148.000 ;
		LAYER M5 ;
		RECT 43.750 146.000 60.445 148.000 ;
		LAYER M5 ;
		RECT 2.000 162.000 27.970 164.000 ;
		LAYER M5 ;
		RECT 43.750 162.000 60.445 164.000 ;

		# Mc2Finalize block inhibit statement blockage
		# Promoted blockages
		LAYER M1 ;
		RECT 57.355 0.000 58.155 0.520 ;
		LAYER M1 ;
		RECT 56.435 0.000 56.515 0.520 ;
		LAYER M2 ;
		RECT 56.435 0.000 56.515 0.520 ;
		LAYER M3 ;
		RECT 56.435 0.000 56.515 0.520 ;
		LAYER M3 ;
		RECT 57.355 0.000 58.155 0.520 ;
		LAYER M2 ;
		RECT 57.355 0.000 58.155 0.520 ;
		LAYER M2 ;
		RECT 58.995 0.000 59.795 0.520 ;
		LAYER M1 ;
		RECT 54.795 0.000 55.595 0.520 ;
		LAYER M2 ;
		RECT 54.795 0.000 55.595 0.520 ;
		LAYER M1 ;
		RECT 58.995 0.000 59.795 0.520 ;
		LAYER M3 ;
		RECT 58.995 0.000 59.795 0.520 ;
		LAYER M3 ;
		RECT 54.795 0.000 55.595 0.520 ;
		LAYER M2 ;
		RECT 60.635 0.000 62.445 0.520 ;
		LAYER M3 ;
		RECT 60.635 0.000 62.445 0.520 ;
		LAYER M1 ;
		RECT 53.155 0.000 53.955 0.520 ;
		LAYER M1 ;
		RECT 60.635 0.000 62.445 0.520 ;
		LAYER M2 ;
		RECT 53.155 0.000 53.955 0.520 ;
		LAYER M3 ;
		RECT 53.155 0.000 53.955 0.520 ;
		LAYER M3 ;
		RECT 41.920 0.000 47.510 0.520 ;
		LAYER M1 ;
		RECT 48.350 0.000 50.565 0.520 ;
		LAYER M3 ;
		RECT 48.350 0.000 50.565 0.520 ;
		LAYER M2 ;
		RECT 48.350 0.000 50.565 0.520 ;
		LAYER M1 ;
		RECT 52.125 0.000 52.315 0.520 ;
		LAYER M3 ;
		RECT 52.125 0.000 52.315 0.520 ;
		LAYER M2 ;
		RECT 52.125 0.000 52.315 0.520 ;
		LAYER M1 ;
		RECT 6.850 0.000 7.650 0.520 ;
		LAYER M2 ;
		RECT 6.850 0.000 7.650 0.520 ;
		LAYER M1 ;
		RECT 16.070 0.000 17.110 0.520 ;
		LAYER M2 ;
		RECT 16.070 0.000 17.110 0.520 ;
		LAYER M3 ;
		RECT 16.070 0.000 17.110 0.520 ;
		LAYER M3 ;
		RECT 6.850 0.000 7.650 0.520 ;
		LAYER M1 ;
		RECT 8.490 0.000 9.290 0.520 ;
		LAYER M2 ;
		RECT 8.490 0.000 9.290 0.520 ;
		LAYER M1 ;
		RECT 10.130 0.000 15.230 0.520 ;
		LAYER M2 ;
		RECT 10.130 0.000 15.230 0.520 ;
		LAYER M3 ;
		RECT 10.130 0.000 15.230 0.520 ;
		LAYER M3 ;
		RECT 8.490 0.000 9.290 0.520 ;
		LAYER M1 ;
		RECT 41.920 0.000 47.510 0.520 ;
		LAYER M2 ;
		RECT 41.920 0.000 47.510 0.520 ;
		LAYER M2 ;
		RECT 36.675 0.000 39.615 0.520 ;
		LAYER M2 ;
		RECT 34.075 0.000 35.835 0.520 ;
		LAYER M2 ;
		RECT 40.455 0.000 41.080 0.520 ;
		LAYER M3 ;
		RECT 36.675 0.000 39.615 0.520 ;
		LAYER M1 ;
		RECT 36.675 0.000 39.615 0.520 ;
		LAYER M1 ;
		RECT 40.455 0.000 41.080 0.520 ;
		LAYER M3 ;
		RECT 40.455 0.000 41.080 0.520 ;
		LAYER M3 ;
		RECT 34.075 0.000 35.835 0.520 ;
		LAYER M1 ;
		RECT 5.930 0.000 6.010 0.520 ;
		LAYER M2 ;
		RECT 5.930 0.000 6.010 0.520 ;
		LAYER M3 ;
		RECT 5.930 0.000 6.010 0.520 ;
		LAYER M4 ;
		RECT 1.415 0.730 1.580 181.555 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 62.445 181.555 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 62.445 181.555 ;
		LAYER M1 ;
		RECT 0.000 0.000 1.810 181.555 ;
		LAYER M2 ;
		RECT 0.000 0.000 1.810 181.555 ;
		LAYER M3 ;
		RECT 0.000 0.000 1.810 181.555 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 62.445 181.555 ;
		LAYER M1 ;
		RECT 17.950 0.000 18.990 0.520 ;
		LAYER M1 ;
		RECT 19.830 0.000 22.750 0.520 ;
		LAYER M2 ;
		RECT 31.110 0.000 32.150 0.520 ;
		LAYER M2 ;
		RECT 19.830 0.000 22.750 0.520 ;
		LAYER M3 ;
		RECT 19.830 0.000 22.750 0.520 ;
		LAYER M3 ;
		RECT 17.950 0.000 18.990 0.520 ;
		LAYER M1 ;
		RECT 23.590 0.000 24.630 0.520 ;
		LAYER M3 ;
		RECT 23.590 0.000 24.630 0.520 ;
		LAYER M3 ;
		RECT 27.350 0.000 30.270 0.520 ;
		LAYER M2 ;
		RECT 23.590 0.000 24.630 0.520 ;
		LAYER M1 ;
		RECT 31.110 0.000 32.150 0.520 ;
		LAYER M2 ;
		RECT 27.350 0.000 30.270 0.520 ;
		LAYER M3 ;
		RECT 31.110 0.000 32.150 0.520 ;
		LAYER M2 ;
		RECT 17.950 0.000 18.990 0.520 ;
		LAYER M1 ;
		RECT 32.990 0.000 33.235 0.520 ;
		LAYER M3 ;
		RECT 32.990 0.000 33.235 0.520 ;
		LAYER M1 ;
		RECT 25.470 0.000 26.510 0.520 ;
		LAYER M2 ;
		RECT 25.470 0.000 26.510 0.520 ;
		LAYER M3 ;
		RECT 25.470 0.000 26.510 0.520 ;
		LAYER M1 ;
		RECT 27.350 0.000 30.270 0.520 ;
		LAYER M3 ;
		RECT 2.650 0.000 3.450 0.520 ;
		LAYER M1 ;
		RECT 2.650 0.000 3.450 0.520 ;
		LAYER M2 ;
		RECT 2.650 0.000 3.450 0.520 ;
		LAYER M4 ;
		RECT 22.310 0.730 22.810 181.555 ;
		LAYER M2 ;
		RECT 32.990 0.000 33.235 0.520 ;
		LAYER M1 ;
		RECT 34.075 0.000 35.835 0.520 ;
		LAYER M4 ;
		RECT 60.865 0.730 61.030 181.555 ;
		LAYER M4 ;
		RECT 49.820 0.730 49.985 181.555 ;
		LAYER M4 ;
		RECT 48.875 0.730 49.440 181.555 ;
		LAYER M1 ;
		RECT 1.810 0.520 62.445 181.555 ;
		LAYER M4 ;
		RECT 10.360 0.730 10.525 181.555 ;
		LAYER M3 ;
		RECT 1.810 0.520 62.445 181.555 ;
		LAYER M2 ;
		RECT 4.290 0.000 5.090 0.520 ;
		LAYER M3 ;
		RECT 4.290 0.000 5.090 0.520 ;
		LAYER M1 ;
		RECT 4.290 0.000 5.090 0.520 ;
		LAYER M2 ;
		RECT 1.810 0.520 62.445 181.555 ;
	END
	# End of OBS

END TS1N65LPA1024X4M4

END LIBRARY

# Created by MC2 : Version 2006.09.01.d on 2024/04/08, 13:51:02

###############################################################################
#        Software       : TSMC MEMORY COMPILER 2006.09.01.d
#        Technology     : 65 nm CMOS LOGIC Low Power LowK Cu 1P9M 1.2
#                         Mix-vt logic, High-vt SRAM
#        Memory Type    : TSMC 65nm low power SP SRAM Without Redundancy
#        Library Name   : ts1n65lpa256x8m4
#        Library Version: 140a
#        Generated Time : 2024/04/08, 13:51:00
###############################################################################
#
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
#
###############################################################################
 
MACRO TS1N65LPA256X8M4
	CLASS BLOCK ;
	FOREIGN TS1N65LPA256X8M4 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 75.965 BY 83.155 ;
	SYMMETRY X Y R90 ;

	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 34.275 0.000 34.795 0.520 ;
			LAYER M1 ;
			RECT 34.275 0.000 34.795 0.520 ;
			LAYER M2 ;
			RECT 34.275 0.000 34.795 0.520 ;
		END
	END A[0]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 36.875 0.000 37.395 0.520 ;
			LAYER M3 ;
			RECT 36.875 0.000 37.395 0.520 ;
			LAYER M1 ;
			RECT 36.875 0.000 37.395 0.520 ;
		END
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 33.190 0.000 33.710 0.520 ;
			LAYER M3 ;
			RECT 33.190 0.000 33.710 0.520 ;
			LAYER M2 ;
			RECT 33.190 0.000 33.710 0.520 ;
		END
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 31.310 0.000 31.830 0.520 ;
			LAYER M3 ;
			RECT 31.310 0.000 31.830 0.520 ;
			LAYER M1 ;
			RECT 31.310 0.000 31.830 0.520 ;
		END
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 27.550 0.000 28.070 0.520 ;
			LAYER M2 ;
			RECT 27.550 0.000 28.070 0.520 ;
			LAYER M1 ;
			RECT 27.550 0.000 28.070 0.520 ;
		END
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 23.120 0.000 23.640 0.520 ;
			LAYER M3 ;
			RECT 23.120 0.000 23.640 0.520 ;
			LAYER M2 ;
			RECT 23.120 0.000 23.640 0.520 ;
		END
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 25.720 0.000 26.240 0.520 ;
			LAYER M1 ;
			RECT 25.720 0.000 26.240 0.520 ;
			LAYER M3 ;
			RECT 25.720 0.000 26.240 0.520 ;
		END
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 19.360 0.000 19.880 0.520 ;
			LAYER M3 ;
			RECT 19.360 0.000 19.880 0.520 ;
			LAYER M1 ;
			RECT 19.360 0.000 19.880 0.520 ;
		END
	END A[7]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 5.250 0.000 5.770 0.520 ;
			LAYER M2 ;
			RECT 5.250 0.000 5.770 0.520 ;
			LAYER M1 ;
			RECT 5.250 0.000 5.770 0.520 ;
		END
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 9.450 0.000 9.970 0.520 ;
			LAYER M1 ;
			RECT 9.450 0.000 9.970 0.520 ;
			LAYER M3 ;
			RECT 9.450 0.000 9.970 0.520 ;
		END
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 13.650 0.000 14.170 0.520 ;
			LAYER M1 ;
			RECT 13.650 0.000 14.170 0.520 ;
			LAYER M3 ;
			RECT 13.650 0.000 14.170 0.520 ;
		END
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 17.850 0.000 18.370 0.520 ;
			LAYER M1 ;
			RECT 17.850 0.000 18.370 0.520 ;
			LAYER M2 ;
			RECT 17.850 0.000 18.370 0.520 ;
		END
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.595 0.000 58.115 0.520 ;
			LAYER M3 ;
			RECT 57.595 0.000 58.115 0.520 ;
			LAYER M2 ;
			RECT 57.595 0.000 58.115 0.520 ;
		END
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 61.795 0.000 62.315 0.520 ;
			LAYER M1 ;
			RECT 61.795 0.000 62.315 0.520 ;
			LAYER M3 ;
			RECT 61.795 0.000 62.315 0.520 ;
		END
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 65.995 0.000 66.515 0.520 ;
			LAYER M1 ;
			RECT 65.995 0.000 66.515 0.520 ;
			LAYER M3 ;
			RECT 65.995 0.000 66.515 0.520 ;
		END
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 70.195 0.000 70.715 0.520 ;
			LAYER M2 ;
			RECT 70.195 0.000 70.715 0.520 ;
			LAYER M3 ;
			RECT 70.195 0.000 70.715 0.520 ;
		END
	END BWEB[7]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 42.120 0.000 42.640 0.520 ;
			LAYER M3 ;
			RECT 42.120 0.000 42.640 0.520 ;
			LAYER M1 ;
			RECT 42.120 0.000 42.640 0.520 ;
		END
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 48.550 0.000 49.070 0.520 ;
			LAYER M1 ;
			RECT 48.550 0.000 49.070 0.520 ;
			LAYER M2 ;
			RECT 48.550 0.000 49.070 0.520 ;
		END
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 1.970 0.000 2.490 0.520 ;
			LAYER M3 ;
			RECT 1.970 0.000 2.490 0.520 ;
			LAYER M1 ;
			RECT 1.970 0.000 2.490 0.520 ;
		END
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 6.170 0.000 6.690 0.520 ;
			LAYER M2 ;
			RECT 6.170 0.000 6.690 0.520 ;
			LAYER M3 ;
			RECT 6.170 0.000 6.690 0.520 ;
		END
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 10.370 0.000 10.890 0.520 ;
			LAYER M1 ;
			RECT 10.370 0.000 10.890 0.520 ;
			LAYER M3 ;
			RECT 10.370 0.000 10.890 0.520 ;
		END
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 14.570 0.000 15.090 0.520 ;
			LAYER M3 ;
			RECT 14.570 0.000 15.090 0.520 ;
			LAYER M1 ;
			RECT 14.570 0.000 15.090 0.520 ;
		END
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 60.875 0.000 61.395 0.520 ;
			LAYER M3 ;
			RECT 60.875 0.000 61.395 0.520 ;
			LAYER M1 ;
			RECT 60.875 0.000 61.395 0.520 ;
		END
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 65.075 0.000 65.595 0.520 ;
			LAYER M3 ;
			RECT 65.075 0.000 65.595 0.520 ;
			LAYER M1 ;
			RECT 65.075 0.000 65.595 0.520 ;
		END
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 69.275 0.000 69.795 0.520 ;
			LAYER M2 ;
			RECT 69.275 0.000 69.795 0.520 ;
			LAYER M3 ;
			RECT 69.275 0.000 69.795 0.520 ;
		END
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 73.475 0.000 73.995 0.520 ;
			LAYER M1 ;
			RECT 73.475 0.000 73.995 0.520 ;
			LAYER M2 ;
			RECT 73.475 0.000 73.995 0.520 ;
		END
	END D[7]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 3.610 0.000 4.130 0.520 ;
			LAYER M1 ;
			RECT 3.610 0.000 4.130 0.520 ;
			LAYER M3 ;
			RECT 3.610 0.000 4.130 0.520 ;
		END
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 7.810 0.000 8.330 0.520 ;
			LAYER M1 ;
			RECT 7.810 0.000 8.330 0.520 ;
			LAYER M3 ;
			RECT 7.810 0.000 8.330 0.520 ;
		END
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 12.010 0.000 12.530 0.520 ;
			LAYER M1 ;
			RECT 12.010 0.000 12.530 0.520 ;
			LAYER M3 ;
			RECT 12.010 0.000 12.530 0.520 ;
		END
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 16.210 0.000 16.730 0.520 ;
			LAYER M1 ;
			RECT 16.210 0.000 16.730 0.520 ;
			LAYER M3 ;
			RECT 16.210 0.000 16.730 0.520 ;
		END
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 59.235 0.000 59.755 0.520 ;
			LAYER M3 ;
			RECT 59.235 0.000 59.755 0.520 ;
			LAYER M1 ;
			RECT 59.235 0.000 59.755 0.520 ;
		END
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 63.435 0.000 63.955 0.520 ;
			LAYER M3 ;
			RECT 63.435 0.000 63.955 0.520 ;
			LAYER M1 ;
			RECT 63.435 0.000 63.955 0.520 ;
		END
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 67.635 0.000 68.155 0.520 ;
			LAYER M3 ;
			RECT 67.635 0.000 68.155 0.520 ;
			LAYER M1 ;
			RECT 67.635 0.000 68.155 0.520 ;
		END
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 71.835 0.000 72.355 0.520 ;
			LAYER M3 ;
			RECT 71.835 0.000 72.355 0.520 ;
			LAYER M1 ;
			RECT 71.835 0.000 72.355 0.520 ;
		END
	END Q[7]

	PIN TSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 52.325 0.000 52.845 0.520 ;
			LAYER M3 ;
			RECT 52.325 0.000 52.845 0.520 ;
			LAYER M1 ;
			RECT 52.325 0.000 52.845 0.520 ;
		END
	END TSEL[0]

	PIN TSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 51.605 0.000 52.125 0.520 ;
			LAYER M3 ;
			RECT 51.605 0.000 52.125 0.520 ;
			LAYER M1 ;
			RECT 51.605 0.000 52.125 0.520 ;
		END
	END TSEL[1]

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 40.655 0.000 41.175 0.520 ;
			LAYER M2 ;
			RECT 40.655 0.000 41.175 0.520 ;
			LAYER M1 ;
			RECT 40.655 0.000 41.175 0.520 ;
		END
	END WEB
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M5 ;
			RECT 0.000 10.000 35.090 14.000 ;
			LAYER M5 ;
			RECT 46.870 10.000 75.965 14.000 ;
			LAYER M5 ;
			RECT 0.000 26.000 35.090 30.000 ;
			LAYER M5 ;
			RECT 46.870 26.000 75.965 30.000 ;
			LAYER M5 ;
			RECT 0.000 42.000 35.090 46.000 ;
			LAYER M5 ;
			RECT 46.870 42.000 75.965 46.000 ;
			LAYER M5 ;
			RECT 0.000 58.000 35.090 62.000 ;
			LAYER M5 ;
			RECT 46.870 58.000 75.965 62.000 ;
			LAYER M5 ;
			RECT 0.000 74.000 35.090 78.000 ;
			LAYER M5 ;
			RECT 46.870 74.000 75.965 78.000 ;
		LAYER M4 ;
		RECT 0.140 0.730 0.470 83.155 ;
		LAYER M4 ;
		RECT 1.580 0.730 1.960 83.155 ;
		LAYER M4 ;
		RECT 3.680 0.730 4.060 83.155 ;
		LAYER M4 ;
		RECT 5.780 0.730 6.160 83.155 ;
		LAYER M4 ;
		RECT 7.880 0.730 8.260 83.155 ;
		LAYER M4 ;
		RECT 9.980 0.730 10.360 83.155 ;
		LAYER M4 ;
		RECT 12.080 0.730 12.460 83.155 ;
		LAYER M4 ;
		RECT 14.180 0.730 14.560 83.155 ;
		LAYER M4 ;
		RECT 16.280 0.730 16.660 83.155 ;
		LAYER M4 ;
		RECT 18.380 0.730 18.760 83.155 ;
		LAYER M4 ;
		RECT 27.930 0.730 30.930 83.155 ;
		LAYER M4 ;
		RECT 39.430 0.730 41.430 83.155 ;
		LAYER M4 ;
		RECT 46.870 0.730 48.870 83.155 ;
		LAYER M4 ;
		RECT 55.105 0.730 55.485 83.155 ;
		LAYER M4 ;
		RECT 57.205 0.730 57.585 83.155 ;
		LAYER M4 ;
		RECT 59.305 0.730 59.685 83.155 ;
		LAYER M4 ;
		RECT 61.405 0.730 61.785 83.155 ;
		LAYER M4 ;
		RECT 63.505 0.730 63.885 83.155 ;
		LAYER M4 ;
		RECT 65.605 0.730 65.985 83.155 ;
		LAYER M4 ;
		RECT 67.705 0.730 68.085 83.155 ;
		LAYER M4 ;
		RECT 69.805 0.730 70.185 83.155 ;
		LAYER M4 ;
		RECT 71.905 0.730 72.285 83.155 ;
		LAYER M4 ;
		RECT 74.005 0.730 74.385 83.155 ;
		LAYER M4 ;
		RECT 75.495 0.730 75.825 83.155 ;
		END
	END VDD

	PIN GND
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M5 ;
			RECT 0.000 2.000 35.090 6.000 ;
			LAYER M5 ;
			RECT 46.870 2.000 75.965 6.000 ;
			LAYER M5 ;
			RECT 0.000 18.000 35.090 22.000 ;
			LAYER M5 ;
			RECT 46.870 18.000 75.965 22.000 ;
			LAYER M5 ;
			RECT 0.000 34.000 35.090 38.000 ;
			LAYER M5 ;
			RECT 46.870 34.000 75.965 38.000 ;
			LAYER M5 ;
			RECT 0.000 50.000 35.090 54.000 ;
			LAYER M5 ;
			RECT 46.870 50.000 75.965 54.000 ;
			LAYER M5 ;
			RECT 0.000 66.000 35.090 70.000 ;
			LAYER M5 ;
			RECT 46.870 66.000 75.965 70.000 ;
		LAYER M4 ;
		RECT 18.925 0.730 19.305 83.155 ;
		LAYER M4 ;
		RECT 27.030 0.730 27.430 83.155 ;
		LAYER M4 ;
		RECT 32.390 0.730 35.090 83.155 ;
		LAYER M4 ;
		RECT 50.795 0.730 53.995 83.155 ;
		LAYER M4 ;
		RECT 54.560 0.730 54.940 83.155 ;
		LAYER M4 ;
		RECT 56.055 0.730 56.635 83.155 ;
		LAYER M4 ;
		RECT 1.035 0.730 1.415 83.155 ;
		LAYER M4 ;
		RECT 2.530 0.730 3.110 83.155 ;
		LAYER M4 ;
		RECT 4.630 0.730 5.210 83.155 ;
		LAYER M4 ;
		RECT 6.730 0.730 7.310 83.155 ;
		LAYER M4 ;
		RECT 8.830 0.730 9.410 83.155 ;
		LAYER M4 ;
		RECT 10.930 0.730 11.510 83.155 ;
		LAYER M4 ;
		RECT 13.030 0.730 13.610 83.155 ;
		LAYER M4 ;
		RECT 15.130 0.730 15.710 83.155 ;
		LAYER M4 ;
		RECT 17.230 0.730 17.810 83.155 ;
		LAYER M4 ;
		RECT 58.155 0.730 58.735 83.155 ;
		LAYER M4 ;
		RECT 60.255 0.730 60.835 83.155 ;
		LAYER M4 ;
		RECT 62.355 0.730 62.935 83.155 ;
		LAYER M4 ;
		RECT 64.455 0.730 65.035 83.155 ;
		LAYER M4 ;
		RECT 66.555 0.730 67.135 83.155 ;
		LAYER M4 ;
		RECT 68.655 0.730 69.235 83.155 ;
		LAYER M4 ;
		RECT 70.755 0.730 71.335 83.155 ;
		LAYER M4 ;
		RECT 72.855 0.730 73.435 83.155 ;
		LAYER M4 ;
		RECT 74.550 0.730 74.930 83.155 ;
		END
	END GND

	OBS
		# Pmesh blockages
		LAYER M5 ;
		RECT 2.000 10.000 33.090 12.000 ;
		LAYER M5 ;
		RECT 48.870 10.000 73.965 12.000 ;
		LAYER M5 ;
		RECT 2.000 26.000 33.090 28.000 ;
		LAYER M5 ;
		RECT 48.870 26.000 73.965 28.000 ;
		LAYER M5 ;
		RECT 2.000 42.000 33.090 44.000 ;
		LAYER M5 ;
		RECT 48.870 42.000 73.965 44.000 ;
		LAYER M5 ;
		RECT 2.000 58.000 33.090 60.000 ;
		LAYER M5 ;
		RECT 48.870 58.000 73.965 60.000 ;
		LAYER M5 ;
		RECT 2.000 74.000 33.090 76.000 ;
		LAYER M5 ;
		RECT 48.870 74.000 73.965 76.000 ;
		LAYER M5 ;
		RECT 2.000 2.000 33.090 4.000 ;
		LAYER M5 ;
		RECT 48.870 2.000 73.965 4.000 ;
		LAYER M5 ;
		RECT 2.000 18.000 33.090 20.000 ;
		LAYER M5 ;
		RECT 48.870 18.000 73.965 20.000 ;
		LAYER M5 ;
		RECT 2.000 34.000 33.090 36.000 ;
		LAYER M5 ;
		RECT 48.870 34.000 73.965 36.000 ;
		LAYER M5 ;
		RECT 2.000 50.000 33.090 52.000 ;
		LAYER M5 ;
		RECT 48.870 50.000 73.965 52.000 ;
		LAYER M5 ;
		RECT 2.000 66.000 33.090 68.000 ;
		LAYER M5 ;
		RECT 48.870 66.000 73.965 68.000 ;

		# Mc2Finalize block inhibit statement blockage
		# Promoted blockages
		LAYER M1 ;
		RECT 70.875 0.000 71.675 0.520 ;
		LAYER M1 ;
		RECT 6.850 0.000 7.650 0.520 ;
		LAYER M3 ;
		RECT 6.850 0.000 7.650 0.520 ;
		LAYER M2 ;
		RECT 6.850 0.000 7.650 0.520 ;
		LAYER M1 ;
		RECT 66.675 0.000 67.475 0.520 ;
		LAYER M3 ;
		RECT 64.115 0.000 64.915 0.520 ;
		LAYER M1 ;
		RECT 64.115 0.000 64.915 0.520 ;
		LAYER M2 ;
		RECT 64.115 0.000 64.915 0.520 ;
		LAYER M2 ;
		RECT 62.475 0.000 63.275 0.520 ;
		LAYER M1 ;
		RECT 62.475 0.000 63.275 0.520 ;
		LAYER M3 ;
		RECT 62.475 0.000 63.275 0.520 ;
		LAYER M2 ;
		RECT 59.915 0.000 60.715 0.520 ;
		LAYER M3 ;
		RECT 59.915 0.000 60.715 0.520 ;
		LAYER M2 ;
		RECT 58.275 0.000 59.075 0.520 ;
		LAYER M1 ;
		RECT 53.005 0.000 57.435 0.520 ;
		LAYER M1 ;
		RECT 58.275 0.000 59.075 0.520 ;
		LAYER M3 ;
		RECT 58.275 0.000 59.075 0.520 ;
		LAYER M2 ;
		RECT 65.755 0.000 65.835 0.520 ;
		LAYER M1 ;
		RECT 61.555 0.000 61.635 0.520 ;
		LAYER M1 ;
		RECT 59.915 0.000 60.715 0.520 ;
		LAYER M2 ;
		RECT 61.555 0.000 61.635 0.520 ;
		LAYER M3 ;
		RECT 61.555 0.000 61.635 0.520 ;
		LAYER M1 ;
		RECT 69.955 0.000 70.035 0.520 ;
		LAYER M2 ;
		RECT 69.955 0.000 70.035 0.520 ;
		LAYER M3 ;
		RECT 69.955 0.000 70.035 0.520 ;
		LAYER M1 ;
		RECT 68.315 0.000 69.115 0.520 ;
		LAYER M2 ;
		RECT 68.315 0.000 69.115 0.520 ;
		LAYER M3 ;
		RECT 68.315 0.000 69.115 0.520 ;
		LAYER M2 ;
		RECT 70.875 0.000 71.675 0.520 ;
		LAYER M3 ;
		RECT 70.875 0.000 71.675 0.520 ;
		LAYER M3 ;
		RECT 72.515 0.000 73.315 0.520 ;
		LAYER M2 ;
		RECT 72.515 0.000 73.315 0.520 ;
		LAYER M1 ;
		RECT 72.515 0.000 73.315 0.520 ;
		LAYER M3 ;
		RECT 66.675 0.000 67.475 0.520 ;
		LAYER M2 ;
		RECT 66.675 0.000 67.475 0.520 ;
		LAYER M3 ;
		RECT 65.755 0.000 65.835 0.520 ;
		LAYER M1 ;
		RECT 65.755 0.000 65.835 0.520 ;
		LAYER M1 ;
		RECT 5.930 0.000 6.010 0.520 ;
		LAYER M3 ;
		RECT 5.930 0.000 6.010 0.520 ;
		LAYER M2 ;
		RECT 5.930 0.000 6.010 0.520 ;
		LAYER M1 ;
		RECT 18.530 0.000 19.200 0.520 ;
		LAYER M3 ;
		RECT 15.250 0.000 16.050 0.520 ;
		LAYER M3 ;
		RECT 20.040 0.000 22.960 0.520 ;
		LAYER M2 ;
		RECT 20.040 0.000 22.960 0.520 ;
		LAYER M1 ;
		RECT 20.040 0.000 22.960 0.520 ;
		LAYER M2 ;
		RECT 18.530 0.000 19.200 0.520 ;
		LAYER M1 ;
		RECT 14.330 0.000 14.410 0.520 ;
		LAYER M1 ;
		RECT 12.690 0.000 13.490 0.520 ;
		LAYER M2 ;
		RECT 12.690 0.000 13.490 0.520 ;
		LAYER M2 ;
		RECT 14.330 0.000 14.410 0.520 ;
		LAYER M3 ;
		RECT 14.330 0.000 14.410 0.520 ;
		LAYER M3 ;
		RECT 18.530 0.000 19.200 0.520 ;
		LAYER M1 ;
		RECT 11.050 0.000 11.850 0.520 ;
		LAYER M3 ;
		RECT 12.690 0.000 13.490 0.520 ;
		LAYER M2 ;
		RECT 11.050 0.000 11.850 0.520 ;
		LAYER M3 ;
		RECT 31.990 0.000 33.030 0.520 ;
		LAYER M1 ;
		RECT 23.800 0.000 25.560 0.520 ;
		LAYER M2 ;
		RECT 26.400 0.000 27.390 0.520 ;
		LAYER M2 ;
		RECT 16.890 0.000 17.690 0.520 ;
		LAYER M1 ;
		RECT 16.890 0.000 17.690 0.520 ;
		LAYER M2 ;
		RECT 15.250 0.000 16.050 0.520 ;
		LAYER M1 ;
		RECT 15.250 0.000 16.050 0.520 ;
		LAYER M2 ;
		RECT 28.230 0.000 31.150 0.520 ;
		LAYER M1 ;
		RECT 28.230 0.000 31.150 0.520 ;
		LAYER M3 ;
		RECT 28.230 0.000 31.150 0.520 ;
		LAYER M1 ;
		RECT 26.400 0.000 27.390 0.520 ;
		LAYER M3 ;
		RECT 26.400 0.000 27.390 0.520 ;
		LAYER M3 ;
		RECT 53.005 0.000 57.435 0.520 ;
		LAYER M2 ;
		RECT 53.005 0.000 57.435 0.520 ;
		LAYER M1 ;
		RECT 49.230 0.000 51.445 0.520 ;
		LAYER M3 ;
		RECT 49.230 0.000 51.445 0.520 ;
		LAYER M2 ;
		RECT 49.230 0.000 51.445 0.520 ;
		LAYER M2 ;
		RECT 42.800 0.000 48.390 0.520 ;
		LAYER M3 ;
		RECT 23.800 0.000 25.560 0.520 ;
		LAYER M2 ;
		RECT 23.800 0.000 25.560 0.520 ;
		LAYER M1 ;
		RECT 42.800 0.000 48.390 0.520 ;
		LAYER M3 ;
		RECT 42.800 0.000 48.390 0.520 ;
		LAYER M1 ;
		RECT 41.335 0.000 41.960 0.520 ;
		LAYER M1 ;
		RECT 37.555 0.000 40.495 0.520 ;
		LAYER M2 ;
		RECT 37.555 0.000 40.495 0.520 ;
		LAYER M2 ;
		RECT 41.335 0.000 41.960 0.520 ;
		LAYER M3 ;
		RECT 41.335 0.000 41.960 0.520 ;
		LAYER M3 ;
		RECT 37.555 0.000 40.495 0.520 ;
		LAYER M3 ;
		RECT 33.870 0.000 34.115 0.520 ;
		LAYER M1 ;
		RECT 33.870 0.000 34.115 0.520 ;
		LAYER M2 ;
		RECT 33.870 0.000 34.115 0.520 ;
		LAYER M1 ;
		RECT 34.955 0.000 36.715 0.520 ;
		LAYER M2 ;
		RECT 34.955 0.000 36.715 0.520 ;
		LAYER M3 ;
		RECT 34.955 0.000 36.715 0.520 ;
		LAYER M2 ;
		RECT 2.650 0.000 3.450 0.520 ;
		LAYER M3 ;
		RECT 2.650 0.000 3.450 0.520 ;
		LAYER M1 ;
		RECT 2.650 0.000 3.450 0.520 ;
		LAYER M4 ;
		RECT 74.385 0.730 74.550 83.155 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 75.965 83.155 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 75.965 83.155 ;
		LAYER M3 ;
		RECT 74.155 0.000 75.965 0.520 ;
		LAYER M2 ;
		RECT 4.290 0.000 5.090 0.520 ;
		LAYER M3 ;
		RECT 4.290 0.000 5.090 0.520 ;
		LAYER M1 ;
		RECT 4.290 0.000 5.090 0.520 ;
		LAYER M1 ;
		RECT 74.155 0.000 75.965 0.520 ;
		LAYER M2 ;
		RECT 74.155 0.000 75.965 0.520 ;
		LAYER M4 ;
		RECT 18.760 0.730 18.925 83.155 ;
		LAYER M3 ;
		RECT 1.810 0.520 75.965 83.155 ;
		LAYER M2 ;
		RECT 1.810 0.520 75.965 83.155 ;
		LAYER M4 ;
		RECT 27.430 0.730 27.930 83.155 ;
		LAYER M4 ;
		RECT 1.415 0.730 1.580 83.155 ;
		LAYER M2 ;
		RECT 0.000 0.000 1.810 83.155 ;
		LAYER M3 ;
		RECT 0.000 0.000 1.810 83.155 ;
		LAYER M1 ;
		RECT 0.000 0.000 1.810 83.155 ;
		LAYER M4 ;
		RECT 53.995 0.730 54.560 83.155 ;
		LAYER M4 ;
		RECT 54.940 0.730 55.105 83.155 ;
		LAYER M1 ;
		RECT 1.810 0.520 75.965 83.155 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 75.965 83.155 ;
		LAYER M3 ;
		RECT 16.890 0.000 17.690 0.520 ;
		LAYER M1 ;
		RECT 31.990 0.000 33.030 0.520 ;
		LAYER M2 ;
		RECT 31.990 0.000 33.030 0.520 ;
		LAYER M3 ;
		RECT 11.050 0.000 11.850 0.520 ;
		LAYER M2 ;
		RECT 8.490 0.000 9.290 0.520 ;
		LAYER M3 ;
		RECT 8.490 0.000 9.290 0.520 ;
		LAYER M2 ;
		RECT 10.130 0.000 10.210 0.520 ;
		LAYER M3 ;
		RECT 10.130 0.000 10.210 0.520 ;
		LAYER M1 ;
		RECT 10.130 0.000 10.210 0.520 ;
		LAYER M1 ;
		RECT 8.490 0.000 9.290 0.520 ;
	END
	# End of OBS

END TS1N65LPA256X8M4

END LIBRARY

**** Created by MC2: Version 2006.09.01.d on 2024/04/08, 13:51:02 

*****************************************************************************
* CDL NETLIST:
* CELL NAME: LEAFCELL
* NETLISTED ON: DEC 15 15:43:47 2005
*****************************************************************************


*****************************************************************************
* GLOBAL NET DECLARATIONS
*****************************************************************************
*.GLOBAL VDD GND


*****************************************************************************
* PIN CONTROL STATEMENT
*****************************************************************************
*.PIN VDD GND


*****************************************************************************
* BIPOLAR DECLARATIONS
*****************************************************************************


*.LDD
*.BIPOLAR 
*.DIOAREA

*.OPTION SCALE=10E-6

*****************************************************************************
* PARAMETER STATEMENT
*****************************************************************************
.PARAM


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRK_DMY                                                            *
* LAST TIME SAVED: OCT 12 13:39:22 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BLTRK_DMY FLOAT TRBL TRWL WL
MN0 BL0_IN NET37 GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NET37 BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 TRBL TRWL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MN3 FLOAT WL NET37 GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 NET37 BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN NET37 VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S1100W8_BLTRK_DMY


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRK_EDG                                                            *
* LAST TIME SAVED: JUN 30 15:24:03 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BLTRK_EDG BL_CONT TRWL
MN0 BL0_IN NET37 GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NET37 BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 BL_CONT TRWL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 NET37 BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN NET37 VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S1100W8_BLTRK_EDG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKDUM                                                               *
* LAST TIME SAVED: OCT 12 13:39:16 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_TRKDUM BL_CONT FLOAT TRBL TIEL WL
XBLTRK FLOAT TRBL TIEL WL S1100W8_BLTRK_DMY
XI14 BL_CONT TIEL S1100W8_BLTRK_EDG
.ENDS S1100W8_TRKDUM


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKDUMX2                                                             *
* LAST TIME SAVED: OCT  4 16:07:09 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_TRKDUMX2 BL_CONT[1] BL_CONT[0] TRBL TIEL WL[1] WL[0]
XI45 BL_CONT[1] NET12 TRBL TIEL WL[1] S1100W8_TRKDUM
XI46 BL_CONT[0] NET12 TRBL TIEL WL[0] S1100W8_TRKDUM
.ENDS S1100W8_TRKDUMX2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRK                                                                *
* LAST TIME SAVED: OCT  4 16:01:28 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BLTRK FLOAT TRBL TRBLB TRWL WL
MN0 BL0_IN TRBLB GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NET42 BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 TRBL TRWL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MN3 FLOAT WL NET42 GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 TRBLB BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN TRBLB VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S1100W8_BLTRK


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRK_EDG2                                                           *
* LAST TIME SAVED: JUN 30 15:51:02 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BLTRK_EDG2 BL_CONT BL0_IN NPD2 PPU1 PPU2 TRWL
MN2 BL_CONT TRWL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MN0 BL0_IN TRWL GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NPD2 TRWL GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MP0 PPU2 TRWL VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 PPU1 TRWL VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S1100W8_BLTRK_EDG2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKNOR                                                               *
* LAST TIME SAVED: OCT  4 16:04:22 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_TRKNOR BL_CONT FLOAT TRBL TIEH TRWL WL
XCELTRK FLOAT TRBL TIEH TRWL WL S1100W8_BLTRK
XI18 BL_CONT NET22 NET23 NET20 NET21 TRWL S1100W8_BLTRK_EDG2
.ENDS S1100W8_TRKNOR


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKNORX2                                                             *
* LAST TIME SAVED: JUL  7 17:14:05 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_TRKNORX2 BL_CONT[1] BL_CONT[0] TRBL TIEH TRWL WL[1] WL[0]
XI52 BL_CONT[1] NET17 TRBL TIEH TRWL WL[1] S1100W8_TRKNOR
XI51 BL_CONT[0] NET17 TRBL TIEH TRWL WL[0] S1100W8_TRKNOR
.ENDS S1100W8_TRKNORX2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRKMIN                                                             *
* LAST TIME SAVED: MAY 17 15:57:20 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BLTRKMIN TRBL TRBLB TRWL WL
MN0 BL0_IN TRWL GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NET41 BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 TRBL TRBL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MN3 TRBLB WL NET41 GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 NET41 BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN TRWL VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S1100W8_BLTRKMIN


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRKMIN_EDG                                                         *
* LAST TIME SAVED: JUL  1 10:37:26 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BLTRKMIN_EDG BL_CONT TRBL TRWL
MN0 BL0_IN TRWL GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 TRWL BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 BL_CONT TRBL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 TRWL BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN TRWL VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S1100W8_BLTRKMIN_EDG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKMIN                                                               *
* LAST TIME SAVED: OCT 12 14:09:32 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_TRKMIN BL_CONT TRBL TIEH TRWL WL
XTRK_VCCMIN TRBL TIEH TRWL WL S1100W8_BLTRKMIN
XI23 BL_CONT TRBL TRWL S1100W8_BLTRKMIN_EDG
.ENDS S1100W8_TRKMIN


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKMINX2                                                             *
* LAST TIME SAVED: OCT 12 14:09:24 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_TRKMINX2 BL_CONT[1] BL_CONT[0] TRBL TIEH TRWL WL[1] WL[0]
XI47 BL_CONT[0] TRBL TIEH TRWL WL[0] S1100W8_TRKMIN
XI46 BL_CONT[1] TRBL TIEH TRWL WL[1] S1100W8_TRKMIN
.ENDS S1100W8_TRKMINX2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SINV_HVTP                                                            *
* LAST TIME SAVED: AUG  3 14:45:00 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_SINV_HVTP Y A LN=0.06U WN=0.15U LP=0.06U WP=0.3U
M1 VDD A Y VDD PCH_HVT W=WP L=LP
M0 Y A GND GND NCH W=WN L=LN
.ENDS S1100W8_SINV_HVTP


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SRAM_TIEH                                                            *
* LAST TIME SAVED: OCT 19 14:27:29 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_SRAM_TIEH Z
XI50 Z NET18 S1100W8_SINV_HVTP LN=0.07U WN=2U LP=0.07U WP=8U
MN0 NET18 NET32 GND GND NCH W=0.15U L=0.07U
MP0 VDD NET32 NET32 VDD PCH W=0.3U L=0.07U
MP1 NET32 NET18 VDD VDD PCH W=0.3U L=0.07U
.ENDS S1100W8_SRAM_TIEH


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SINV                                                                 *
* LAST TIME SAVED: APR 15 08:08:15 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_SINV Y A LP=0.06U WP=0.3U LN=0.06U WN=0.15U
M0 Y A GND GND NCH W=WN L=LN
M1 VDD A Y VDD PCH W=WP L=LP
.ENDS S1100W8_SINV


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SNAND3                                                               *
* LAST TIME SAVED: APR 18 16:13:20 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_SNAND3 Y A B C LP3=0.06U WP3=0.3U LP2=0.06U WP2=0.3U LP1=0.06U WP1=0.3U
+LN1=0.06U WN1=0.45U LN2=0.06U WN2=0.45U LN3=0.06U WN3=0.45U
M0 NET14 C GND GND NCH W=WN3 L=LN3
M1 NET17 B NET14 GND NCH W=WN2 L=LN2
M2 Y A NET17 GND NCH W=WN1 L=LN1
M3 VDD A Y VDD PCH W=WP1 L=LP1
M4 VDD B Y VDD PCH W=WP2 L=LP2
M5 VDD C Y VDD PCH W=WP3 L=LP3
.ENDS S1100W8_SNAND3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XDRV                                                                 *
* LAST TIME SAVED: DEC 14 16:50:11 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_XDRV WLOUT[1] WLOUT[0] WLPY WLPYB0 WLPYB1 XPD0 XPD0B XPD1 XPD2
XI288 MWL1 MWL0 S1100W8_SINV LP=0.06U WP=0.8U  LN=0.06U WN=0.8U 
XI295 MWL1A MWL0A S1100W8_SINV LP=0.06U WP=0.8U  LN=0.06U WN=0.8U 
XI296 WLOUT[1] MWL2A S1100W8_SINV_HVTP LN=0.06U WN=5U    LP=0.06U WP=10U    M=2
XI275 WLOUT[0] MWL2 S1100W8_SINV_HVTP LN=0.06U WN=5U    LP=0.06U WP=10U    M=2
MN0 MWL2 MWL1 WLPY GND NCH W=2.0U   L=0.06U
MN1 MWL2A MWL1A WLPY GND NCH W=2.0U   L=0.06U
MP0 VDD MWL1 MWL2 VDD PCH W=2.0U   L=0.06U
MP2 VDD MWL1A MWL2A VDD PCH W=2.0U   L=0.06U
MP3 MWL2A WLPYB0 VDD VDD PCH W=2.0U      L=0.06U
MP1 MWL2 WLPYB1 VDD VDD PCH W=2.0U      L=0.06U
XI290 MWL0A XPD2 XPD1 XPD0B S1100W8_SNAND3 LP3=0.06U WP3=0.15U  LP2=0.06U WP2=0.15U
+LP1=0.06U WP1=0.15U  LN1=0.06U WN1=0.15U  LN2=0.06U WN2=0.15U LN3=0.06U
+WN3=0.15U 
XI282 MWL0 XPD2 XPD1 XPD0 S1100W8_SNAND3 LP3=0.06U WP3=0.15U  LP2=0.06U WP2=0.15U
+LP1=0.06U WP1=0.15U  LN1=0.06U WN1=0.15U  LN2=0.06U WN2=0.15U LN3=0.06U
+WN3=0.15U 
**C2 MWL2 GND 10.372F
**C4 MWL1 GND 3.209F
**C3 MWL0 GND 2.040F
**C5 MWL2A GND 9.991F
**C6 MWL1A GND 3.359F
**C7 MWL0A GND 2.282F
.ENDS S1100W8_XDRV


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XDRVX2                                                               *
* LAST TIME SAVED: JUN 13 11:08:29 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_XDRVX2 WL[3] WL[2] WL[1] WL[0] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2]
+XPD0[1] XPD0[0] XPD1 XPD2
XWLDRV_0 WL[1] WL[0] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1 XPD2 S1100W8_XDRV
XWLDRV_1 WL[2] WL[3] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1 XPD2 S1100W8_XDRV
.ENDS S1100W8_XDRVX2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IOYPASS_M16                                                          *
* LAST TIME SAVED: OCT 12 14:13:51 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IOYPASS_M16 BL BLB DL DLB BLEQB YSEL
*MN0 BL YSEL DL GND NCH W=0.8U L=0.06U
MN0 BL YSEL DL GND NCH W=0.89U L=0.06U
*MN1 BLB YSEL DLB GND NCH W=0.8U L=0.06U
MN1 BLB YSEL DLB GND NCH W=0.89U L=0.06U
MP2 BLB BLEQB BL VDD PCH W=2U L=0.06U
MP0 BL NET47 DL VDD PCH W=0.8U L=0.06U
MP3 VDD BLEQB BLB VDD PCH W=2U L=0.06U
MP1 BLB NET47 DLB VDD PCH W=0.8U L=0.06U
MP4 BL BLEQB VDD VDD PCH W=2U L=0.06U
XI9 NET47 YSEL S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.24U
.ENDS S1100W8_IOYPASS_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DIN                                                                  *
* LAST TIME SAVED: DEC 14 16:50:06 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_DIN AWTD BWEB_M D_M BIST BWEB BWEBM D DM
XI13 BIST_BB BIST_B S1100W8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI12 BIST_B BIST S1100W8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI293 BWEB_M NET16 S1100W8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
XI344 BWC BWT S1100W8_SINV LP=0.15U WP=0.28U LN=0.15U WN=0.15U
XI241 NET14 BWC S1100W8_SINV LP=0.15U WP=0.28U LN=0.15U WN=0.15U
XI242 NET16 NET14 S1100W8_SINV LP=0.1U WP=0.28U LN=0.1U WN=0.15U
XI343 BWT NET107 S1100W8_SINV LP=0.15U WP=0.28U LN=0.15U WN=0.15U
XI85 DT NET110 S1100W8_SINV LP=0.1U WP=0.3U LN=0.1U WN=0.15U
XI83 DC DT S1100W8_SINV LP=0.1U WP=0.3U LN=0.1U WN=0.15U
XI59 D_M NET26 S1100W8_SINV LP=0.07U WP=1.2U LN=0.07U WN=0.6U
XI84 NET26 DC S1100W8_SINV LP=0.2U WP=0.6U LN=0.2U WN=0.3U
**C11 BIST_BB GND 1.596F
**C13 BIST_B GND 1.310F
**C37 NET14 GND 0.680F
**C53 NET16 GND 0.860F
**C23 BWC GND 1.411F
**C14 BWT GND 1.879F
**C12 NET107 GND 1.155F
**C9 DT GND 2.044F
**C2 NET26 GND 1.135F
**C1 DC GND 1.509F
**C10 NET110 GND 1.392F
MP9 NET51 DC AWTD VDD PCH W=0.42U L=0.07U
MP8 VDD BWT NET51 VDD PCH W=0.42U L=0.07U
MP5 VDD BWC NET59 VDD PCH W=0.42U L=0.07U
MP4 NET59 DT AWTD VDD PCH W=0.42U L=0.07U
MP3 NET62 BIST_B NET107 VDD PCH W=0.3U L=0.06U
MP7 VDD BWEBM NET62 VDD PCH W=0.3U L=0.06U
MP1 VDD BWEB NET71 VDD PCH W=0.3U L=0.06U
MP0 NET71 BIST_BB NET107 VDD PCH W=0.3U L=0.06U
MP15 NET74 BIST_BB NET110 VDD PCH W=0.3U L=0.06U
MP14 VDD D NET74 VDD PCH W=0.3U L=0.06U
MP2 VDD DM NET83 VDD PCH W=0.3U L=0.06U
MP6 NET83 BIST_B NET110 VDD PCH W=0.3U L=0.06U
MN7 NET86 BWT GND GND NCH W=0.21U L=0.07U
MN5 AWTD BWC NET86 GND NCH W=0.21U L=0.07U
MN4 AWTD DT NET86 GND NCH W=0.21U L=0.07U
MN3 NET86 DC GND GND NCH W=0.21U L=0.07U
MN6 NET98 BWEBM GND GND NCH W=0.15U L=0.06U
MN2 NET101 BWEB GND GND NCH W=0.15U L=0.06U
MN1 NET107 BIST_BB NET98 GND NCH W=0.15U L=0.06U
MN0 NET107 BIST_B NET101 GND NCH W=0.15U L=0.06U
MN15 NET110 BIST_B NET116 GND NCH W=0.15U L=0.06U
MN14 NET110 BIST_BB NET119 GND NCH W=0.15U L=0.06U
MN13 NET116 D GND GND NCH W=0.15U L=0.06U
MN9 NET119 DM GND GND NCH W=0.15U L=0.06U
.ENDS S1100W8_DIN


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SNOR                                                                 *
* LAST TIME SAVED: APR 15 09:10:54 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_SNOR Y A B LP1=0.06U WP1=0.6U LP2=0.06U WP2=0.6U LN2=0.06U WN2=0.15U LN1=0.06U
+WN1=0.15U
M3 Y A GND GND NCH W=WN1 L=LN1
M2 Y B GND GND NCH W=WN2 L=LN2
M1 NET3 B Y VDD PCH W=WP2 L=LP2
M0 VDD A NET3 VDD PCH W=WP1 L=LP1
.ENDS S1100W8_SNOR


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SA                                                                   *
* LAST TIME SAVED: DEC 14 16:50:07 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_SA Q AWTD AWTI DL DLB PGB PREB SAE
MN11 Z4 AWTD GND GND NCH W=0.9U L=0.07U M=1
MN10 Z4 AWTT Q_B GND NCH W=0.9U L=0.07U M=1
MN8 Z6 AWTC Q_B GND NCH W=0.9U L=0.07U M=1
MN5 Z6 SOB GND GND NCH W=0.9U L=0.07U M=1
MN2 NS SAE GND GND NCH W=2.0U L=0.08U
MN1 DLB_IN DL_IN NS GND NCH W=2.0U L=0.18U
MN0 NS DLB_IN DL_IN GND NCH W=2.0U L=0.18U
MP14 Q_B AWTT Z5 VDD PCH W=1.8U L=0.07U M=1
MP5 Z3 AWTD VDD VDD PCH W=1.8U L=0.07U M=1
MP9 Q_B AWTC Z3 VDD PCH W=1.8U L=0.07U M=1
MP13 Z5 SOB VDD VDD PCH W=1.8U L=0.07U M=1
MP10 VDD PREB DL_IN VDD PCH W=1.0U L=0.1U
MP11 VDD PREB DLB_IN VDD PCH W=1.0U L=0.1U
MP8 DLB_IN PREB DL_IN VDD PCH W=1.2U L=0.12U
MP3 VDD DL_IN DLB_IN VDD PCH W=1.0U L=0.12U
MP2 DL_IN DLB_IN VDD VDD PCH W=1.0U L=0.12U
MP7 DLB PGB DLB_IN VDD PCH W=1.2U L=0.1U
MP6 DL_IN PGB DL VDD PCH W=1.2U L=0.1U
XI152 SO SOB NET096 S1100W8_SNOR LP1=0.07U WP1=2.4U LP2=0.07U WP2=2.4U LN2=0.07U WN2=0.8U
+LN1=0.07U WN1=0.8U
XI116 SOB SO NET098 S1100W8_SNOR LP1=0.07U WP1=2.4U LP2=0.07U WP2=2.4U LN2=0.07U WN2=0.8U
+LN1=0.07U WN1=0.8U
XI153 NET096 DL_IN S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.38U
XI148 NET098 DLB_IN S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.38U
XI61 AWTC AWTI S1100W8_SINV LP=0.06U WP=0.48U LN=0.06U WN=0.24U
XI62 AWTT AWTC S1100W8_SINV LP=0.06U WP=0.48U LN=0.06U WN=0.24U
XI160 Q Q_B S1100W8_SINV LP=0.07U WP=3.6U LN=0.07U WN=1.8U
**C0 DL_IN GND 4.360F
**C1 DLB_IN GND 4.037F
**C4 SO GND 1.951F
**C15 AWTC GND 1.969F
**C7 NET096 GND 2.576F
**C16 AWTT GND 2.078F
**C9 NET098 GND 2.471F
**C14 SOB GND 3.090F
**C17 Q_B GND 2.798F
.ENDS S1100W8_SA


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRANSGATE                                                            *
* LAST TIME SAVED: APR 15 08:43:26 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_TRANSGATE Y A C CB LP=0.06U WP=0.3U LN=0.06U WN=0.15U
*.NOPIN VDD GND
M1 A C Y GND NCH W=WN L=LN
M0 Y CB A VDD PCH W=WP L=LP
.ENDS S1100W8_TRANSGATE


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_DCLK                                                              *
* LAST TIME SAVED: DEC 14 16:50:06 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_LH_DCLK Q CP D
**C2 P2 GND 1.709F
**C0 INCP GND 1.251F
XI26 D P2 CP INCP S1100W8_TRANSGATE LP=0.07U WP=0.5U LN=0.07U WN=0.5U
XI33 Q P2 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI29 INCP CP S1100W8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.3U
MN12 GND Q NET39 GND NCH W=0.15U L=0.07U
MN11 NET39 INCP P2 GND NCH W=0.15U L=0.07U
MP4 NET69 Q VDD VDD PCH W=0.28U L=0.07U
MP5 P2 CP NET69 VDD PCH W=0.28U L=0.07U
.ENDS S1100W8_LH_DCLK


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_WRIN_M16                                                          *
* LAST TIME SAVED: SEP 28 10:50:28 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IO_WRIN_M16 DL DLB D DCLK DLEQB WPG
XLH_DCLK_M8 D1B DCLK D S1100W8_LH_DCLK
MP7 DL DLEQB VDD VDD PCH W=1U L=0.07U
MP8 VDD DLEQB DLB VDD PCH W=1U L=0.07U
MN2 VDD D1 D2B VDD PCH W=2.5U L=0.07U
MN0 VDD D1B D2 VDD PCH W=2.5U L=0.07U
MN5 DLB WPG D2B GND NCH W=2.5U L=0.07U
MN4 D2 WPG DL GND NCH W=2.5U L=0.07U
MN3 D2B D1 GND GND NCH W=5U L=0.07U
MN1 D2 D1B GND GND NCH W=5U L=0.07U
XI69 D1 D1B S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
**C11 D1B GND 4.2F
**C6 D1 GND 2.6F
**C7 D2B GND 4.5F
**C8 D2 GND 4.5F
.ENDS S1100W8_IO_WRIN_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_BWEB                                                              *
* LAST TIME SAVED: DEC 14 16:50:07 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_LH_BWEB Q CP D
MP5 P2 CP NET42 VDD PCH W=0.2U L=0.07U
MP4 NET42 Q VDD VDD PCH W=0.2U L=0.07U
XI26 D P2 CP INCP S1100W8_TRANSGATE LP=0.07U WP=0.5U LN=0.07U WN=0.5U
XI29 INCP CP S1100W8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.2U
XI24 Q P2 S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.4U
MN12 GND Q NET51 GND NCH W=0.2U L=0.07U
MN11 NET51 INCP P2 GND NCH W=0.2U L=0.07U
**C1 P2 GND 1.855F
**C0 INCP GND 1.980F
.ENDS S1100W8_LH_BWEB


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SNAND                                                                *
* LAST TIME SAVED: APR 15 08:59:39 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_SNAND Y A B LP2=0.06U WP2=0.3U LP1=0.06U WP1=0.3U LN1=0.06U WN1=0.3U LN2=0.06U
+WN2=0.3U
M0 NET9 B GND GND NCH W=WN2 L=LN2
M1 Y A NET9 GND NCH W=WN1 L=LN1
M2 VDD A Y VDD PCH W=WP1 L=LP1
M3 VDD B Y VDD PCH W=WP2 L=LP2
.ENDS S1100W8_SNAND


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_RWCTRL_M16                                                        *
* LAST TIME SAVED: OCT  7 14:27:13 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IO_RWCTRL_M16 BLEQB DLEQB DLH PGB PREB SAE WPG BWEB DCLK GW_RB WLP
X_LH_BWEB BWEB_SU DLH BWEB S1100W8_LH_BWEB
XI289 PREB NET0100 NET161 S1100W8_SNOR LP1=0.07U WP1=1.2U LP2=0.07U WP2=1.2U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI288 NET161 WLPCD2 NET163 S1100W8_SNOR LP1=0.07U WP1=0.35U LP2=0.07U WP2=0.35U LN2=0.07U
+WN2=0.3U LN1=0.07U WN1=0.3U
XI249 WPG GW_R NET089 S1100W8_SNOR LP1=0.07U WP1=1.0U LP2=0.07U WP2=1.0U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI133 NET073 WLPCD0 NET_110 GW_R S1100W8_SNAND3 LP3=0.07U WP3=1.75U LP2=0.07U WP2=1.75U
+LP1=0.07U WP1=1.75U LN1=0.07U WN1=1.2U LN2=0.07U WN2=1.2U LN3=0.07U WN3=1.2U
XI250 PGB NET166 GW_R S1100W8_SNAND LP2=0.07U WP2=0.84U LP1=0.07U WP1=0.84U LN1=0.07U
+WN1=0.7U LN2=0.07U WN2=0.7U
XI305 NET90 NET073 WLPCD2 S1100W8_SNAND LP2=0.07U WP2=0.42U LP1=0.07U WP1=0.42U LN1=0.07U
+WN1=0.21U LN2=0.07U WN2=0.21U
XI307 BLEQB WLPCD0 WLPCD4 S1100W8_SNAND LP2=0.07U WP2=1.75U LP1=0.07U WP1=3.5U LN1=0.07U
+WN1=4U LN2=0.07U WN2=4U
XI306 NET289 WLPCD1 BWEB_SU S1100W8_SNAND LP2=0.07U WP2=0.3U LP1=0.07U WP1=0.3U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI339 NET0219 DCLK WLPCD3 S1100W8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI186 NET163 NET93 NET073 S1100W8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI312 NET083 WLPCD0 S1100W8_SINV LP=0.10U WP=0.35U LN=0.10U WN=0.15U
XI73 GW_R GW_RB S1100W8_SINV LP=0.07U WP=1.4U LN=0.07U WN=0.7U
XI348 NET0100 GW_R S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI329 NET0153 WLPCD3 S1100W8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.15U
XI217 WLPCD1 WLPCD0 S1100W8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.28U
XI340 DLH NET0219 S1100W8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.7U
XI287 NET93 NET135 S1100W8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI327 NET141 NET139 S1100W8_SINV LP=0.18U WP=0.35U LN=0.18U WN=0.15U
XI286 NET135 PGB S1100W8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI134 SAE NET073 S1100W8_SINV LP=0.15U WP=0.7U LN=0.1U WN=0.35U
XI321 NET062 NET289 S1100W8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI264 WLPCD4 NET0153 S1100W8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI322 NET089 NET062 S1100W8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.2U
XI185 NET166 NET90 S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.28U
XI299 WLPCD2 NET100 S1100W8_SINV LP=0.07U WP=0.9U LN=0.07U WN=0.3U
XI298 NET100 WLPCD1 S1100W8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI207 NET_110 NET141 S1100W8_SINV LP=0.10U WP=0.7U LN=0.10U WN=0.28U
XI334 DLEQB NET095 S1100W8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
XI337 WLPCD3 WLPCD2 S1100W8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.25U
XI128 WLPCD0 NET085 S1100W8_SINV LP=0.07U WP=1.6U LN=0.07U WN=0.8U
XI315 NET085 WLP S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI333 NET095 BLEQB S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI311 NET088 NET083 S1100W8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
XI310 NET139 NET088 S1100W8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
**C50 WLPCD4 GND 2.8F
**C51 NET135 GND 0.45F
**C17 WLPCD1 GND 1.92F
**C33 NET139 GND 1F
**C15 NET0100 GND 0.57F
**C31 NET_110 GND 2.8F
**C13 NET073 GND 2.95F
**C10 NET095 GND 1.2F
**C11 NET0219 GND 1F
**C48 WLPCD2 GND 2.96F
**C47 NET166 GND 1F
**C26 BWEB_SU GND 1.6F
**C42 NET161 GND 2.1F
**C27 NET93 GND 1.6F
**C43 NET163 GND 0.85F
**C24 NET062 GND 0.7F
**C9 NET0153 GND 0.5F
**C8 WLPCD3 GND 1F
**C7 NET100 GND 0.55F
**C6 NET085 GND 0.6F
**C5 NET089 GND 2.4F
**C4 GW_R GND 4.29F
**C3 NET289 GND 1.1F
**C2 NET083 GND 0.5F
**C1 NET088 GND 1.1F
**C0 NET141 GND 0.7F
**C54 NET90 GND 0.45F
**C18 WLPCD0 GND 4F
.ENDS S1100W8_IO_RWCTRL_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IORWBLK_M16                                                          *
* LAST TIME SAVED: NOV 30 14:33:22 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IORWBLK_M16 BLEQB Q DL DLB AWTI BIST BWEB BWEBM D DCLK DM GW_RB WLP
XDIN AWTD BWEB_M NET46 BIST BWEB BWEBM D DM S1100W8_DIN
XSA Q AWTD AWTI DL DLB PGB PREB SAE S1100W8_SA
XIO_WRIN DL DLB NET46 DCLK_DATA NET041 WPG S1100W8_IO_WRIN_M16
XIO_RWCTRL BLEQB NET041 DCLK_DATA PGB PREB SAE WPG BWEB_M DCLK GW_RB WLP
+S1100W8_IO_RWCTRL_M16
**C3 WPG GND 5F
**C2 SAE GND 5F
**C8 NET041 GND 3.5F
**C4 PGB GND 5F
**C0 DCLK_DATA GND 2F
**C5 PREB GND 5F
**C6 BWEB_M GND 1.7F
**C7 AWTD GND 1.7F
**C1 NET46 GND 1.7F
.ENDS S1100W8_IORWBLK_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YSELX4                                                               *
* LAST TIME SAVED: DEC 12 10:42:39 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_YSELX4 YSEL[3] YSEL[2] YSEL[1] YSEL[0] Y10[3] Y10[2] Y10[1] Y10[0] Y432
**C76 NET15 GND 1.1F
**C77 NET26 GND 1.1F
**C79 NET43 GND 1.1F
**C81 NET40 GND 1.1F
XI73 YSEL[2] NET43 S1100W8_SINV LP=0.07U WP=0.84U LN=0.07U WN=0.41U
XI72 YSEL[1] NET26 S1100W8_SINV LP=0.07U WP=0.84U LN=0.07U WN=0.41U
XI61 YSEL[0] NET15 S1100W8_SINV LP=0.07U WP=0.84U LN=0.07U WN=0.41U
XI74 YSEL[3] NET40 S1100W8_SINV LP=0.07U WP=0.84U LN=0.07U WN=0.41U
MN4 NET40 Y10[3] NET12 GND NCH W=0.32U L=0.07U
MN1 NET15 Y10[0] NET12 GND NCH W=0.32U L=0.07U
MN3 NET43 Y10[2] NET12 GND NCH W=0.32U L=0.07U
MN0 NET12 Y432 GND GND NCH W=0.32U L=0.07U
MN2 NET26 Y10[1] NET12 GND NCH W=0.32U L=0.07U
MP6 VDD Y10[3] NET40 VDD PCH W=0.32U L=0.07U
MP7 VDD Y432 NET40 VDD PCH W=0.32U L=0.07U
MP5 VDD Y432 NET43 VDD PCH W=0.32U L=0.07U
MP3 VDD Y432 NET26 VDD PCH W=0.32U L=0.07U
MP4 VDD Y10[2] NET43 VDD PCH W=0.32U L=0.07U
MP1 VDD Y432 NET15 VDD PCH W=0.32U L=0.07U
MP2 VDD Y10[1] NET26 VDD PCH W=0.32U L=0.07U
MP0 VDD Y10[0] NET15 VDD PCH W=0.32U L=0.07U
.ENDS S1100W8_YSELX4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_M16                                                               *
* LAST TIME SAVED: NOV 10 11:38:59 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IO_M16 Q BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8]
+BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] BLB[2] BLB[3]
+BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14]
+BLB[15] AWTI BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP Y10[3] Y10[2] Y10[1]
+Y10[0] Y32[3] Y32[2] Y32[1] Y32[0]
XIYPASS_15 BL[15] BLB[15] NET25 NET24 NET23 YSEL[15] S1100W8_IOYPASS_M16
XIYPASS_14 BL[14] BLB[14] NET25 NET24 NET23 YSEL[14] S1100W8_IOYPASS_M16
XIYPASS_13 BL[13] BLB[13] NET25 NET24 NET23 YSEL[13] S1100W8_IOYPASS_M16
XIYPASS_12 BL[12] BLB[12] NET25 NET24 NET23 YSEL[12] S1100W8_IOYPASS_M16
XIYPASS_11 BL[11] BLB[11] NET25 NET24 NET23 YSEL[11] S1100W8_IOYPASS_M16
XIYPASS_10 BL[10] BLB[10] NET25 NET24 NET23 YSEL[10] S1100W8_IOYPASS_M16
XIYPASS_9 BL[9] BLB[9] NET25 NET24 NET23 YSEL[9] S1100W8_IOYPASS_M16
XIYPASS_8 BL[8] BLB[8] NET25 NET24 NET23 YSEL[8] S1100W8_IOYPASS_M16
XIYPASS_7 BL[7] BLB[7] NET25 NET24 NET23 YSEL[7] S1100W8_IOYPASS_M16
XIYPASS_6 BL[6] BLB[6] NET25 NET24 NET23 YSEL[6] S1100W8_IOYPASS_M16
XIYPASS_5 BL[5] BLB[5] NET25 NET24 NET23 YSEL[5] S1100W8_IOYPASS_M16
XIYPASS_4 BL[4] BLB[4] NET25 NET24 NET23 YSEL[4] S1100W8_IOYPASS_M16
XIYPASS_3 BL[3] BLB[3] NET25 NET24 NET23 YSEL[3] S1100W8_IOYPASS_M16
XIYPASS_2 BL[2] BLB[2] NET25 NET24 NET23 YSEL[2] S1100W8_IOYPASS_M16
XIYPASS_1 BL[1] BLB[1] NET25 NET24 NET23 YSEL[1] S1100W8_IOYPASS_M16
XIYPASS_0 BL[0] BLB[0] NET25 NET24 NET23 YSEL[0] S1100W8_IOYPASS_M16
XI2 NET23 Q NET25 NET24 AWTI BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP
+S1100W8_IORWBLK_M16
XYSELX4_3 YSEL[15] YSEL[14] YSEL[13] YSEL[12] Y10[3] Y10[2] Y10[1] Y10[0]
+Y32[3] S1100W8_YSELX4
XYSELX4_2 YSEL[11] YSEL[10] YSEL[9] YSEL[8] Y10[3] Y10[2] Y10[1] Y10[0] Y32[2]
+S1100W8_YSELX4
XYSELX4_1 YSEL[7] YSEL[6] YSEL[5] YSEL[4] Y10[3] Y10[2] Y10[1] Y10[0] Y32[1]
+S1100W8_YSELX4
XYSELX4_0 YSEL[3] YSEL[2] YSEL[1] YSEL[0] Y10[3] Y10[2] Y10[1] Y10[0] Y32[0]
+S1100W8_YSELX4
.ENDS S1100W8_IO_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_WRIN_M8                                                           *
* LAST TIME SAVED: SEP 28 10:50:28 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IO_WRIN_M8 DL DLB D DCLK DLEQB WPG
XLH_DCLK_M8 D1B DCLK D S1100W8_LH_DCLK
MP7 DL DLEQB VDD VDD PCH W=1U L=0.07U
MP8 VDD DLEQB DLB VDD PCH W=1U L=0.07U
MN2 VDD D1 D2B VDD PCH W=2.5U L=0.07U
MN0 VDD D1B D2 VDD PCH W=2.5U L=0.07U
MN5 DLB WPG D2B GND NCH W=2.5U L=0.07U
MN4 D2 WPG DL GND NCH W=2.5U L=0.07U
MN3 D2B D1 GND GND NCH W=5U L=0.07U
MN1 D2 D1B GND GND NCH W=5U L=0.07U
XI69 D1 D1B S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
**C11 D1B GND 4.2F
**C6 D1 GND 2.6F
**C7 D2B GND 4.5F
**C8 D2 GND 4.5F
.ENDS S1100W8_IO_WRIN_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_RWCTRL_M8                                                         *
* LAST TIME SAVED: OCT  6 16:44:21 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IO_RWCTRL_M8 BLEQB DLEQB DLH PGB PREB SAE WPG BWEB DCLK GW_RB WLP
X_LH_BWEB BWEB_SU DLH BWEB S1100W8_LH_BWEB
XI289 PREB NET0100 NET161 S1100W8_SNOR LP1=0.07U WP1=1.2U LP2=0.07U WP2=1.2U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI288 NET161 WLPCD2 NET163 S1100W8_SNOR LP1=0.07U WP1=0.35U LP2=0.07U WP2=0.35U LN2=0.07U
+WN2=0.3U LN1=0.07U WN1=0.3U
XI249 WPG GW_R NET089 S1100W8_SNOR LP1=0.07U WP1=1.0U LP2=0.07U WP2=1.0U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI133 NET073 WLPCD0 NET_110 GW_R S1100W8_SNAND3 LP3=0.07U WP3=1.75U LP2=0.07U WP2=1.75U
+LP1=0.07U WP1=1.75U LN1=0.07U WN1=1.2U LN2=0.07U WN2=1.2U LN3=0.07U WN3=1.2U
XI250 PGB NET166 GW_R S1100W8_SNAND LP2=0.07U WP2=0.84U LP1=0.07U WP1=0.84U LN1=0.07U
+WN1=0.7U LN2=0.07U WN2=0.7U
XI305 NET90 NET073 WLPCD2 S1100W8_SNAND LP2=0.07U WP2=0.42U LP1=0.07U WP1=0.42U LN1=0.07U
+WN1=0.21U LN2=0.07U WN2=0.21U
XI307 BLEQB WLPCD0 WLPCD4 S1100W8_SNAND LP2=0.07U WP2=1.75U LP1=0.07U WP1=3.5U LN1=0.07U
+WN1=4U LN2=0.07U WN2=4U
XI306 NET289 WLPCD1 BWEB_SU S1100W8_SNAND LP2=0.07U WP2=0.3U LP1=0.07U WP1=0.3U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI339 NET0219 DCLK WLPCD3 S1100W8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI186 NET163 NET93 NET073 S1100W8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI312 NET083 WLPCD0 S1100W8_SINV LP=0.10U WP=0.35U LN=0.10U WN=0.15U
XI73 GW_R GW_RB S1100W8_SINV LP=0.07U WP=1.4U LN=0.07U WN=0.7U
XI348 NET0100 GW_R S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI329 NET0153 WLPCD3 S1100W8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.15U
XI217 WLPCD1 WLPCD0 S1100W8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.28U
XI340 DLH NET0219 S1100W8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.7U
XI287 NET93 NET135 S1100W8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI327 NET141 NET139 S1100W8_SINV LP=0.18U WP=0.35U LN=0.18U WN=0.15U
XI286 NET135 PGB S1100W8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI134 SAE NET073 S1100W8_SINV LP=0.15U WP=0.7U LN=0.1U WN=0.35U
XI321 NET062 NET289 S1100W8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI264 WLPCD4 NET0153 S1100W8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI322 NET089 NET062 S1100W8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.2U
XI185 NET166 NET90 S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.28U
XI299 WLPCD2 NET100 S1100W8_SINV LP=0.07U WP=0.9U LN=0.07U WN=0.3U
XI298 NET100 WLPCD1 S1100W8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI207 NET_110 NET141 S1100W8_SINV LP=0.10U WP=0.7U LN=0.10U WN=0.28U
XI334 DLEQB NET095 S1100W8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
XI337 WLPCD3 WLPCD2 S1100W8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.25U
XI128 WLPCD0 NET085 S1100W8_SINV LP=0.07U WP=1.6U LN=0.07U WN=0.8U
XI315 NET085 WLP S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI333 NET095 BLEQB S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI311 NET088 NET083 S1100W8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
XI310 NET139 NET088 S1100W8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
**C50 WLPCD4 GND 2.8F
**C51 NET135 GND 0.45F
**C17 WLPCD1 GND 1.92F
**C33 NET139 GND 1F
**C15 NET0100 GND 0.57F
**C31 NET_110 GND 2.8F
**C13 NET073 GND 2.95F
**C10 NET095 GND 1.2F
**C11 NET0219 GND 1F
**C48 WLPCD2 GND 2.96F
**C47 NET166 GND 1F
**C26 BWEB_SU GND 1.6F
**C42 NET161 GND 2.1F
**C27 NET93 GND 1.6F
**C43 NET163 GND 0.85F
**C24 NET062 GND 0.7F
**C9 NET0153 GND 0.5F
**C8 WLPCD3 GND 1F
**C7 NET100 GND 0.55F
**C6 NET085 GND 0.6F
**C5 NET089 GND 2.4F
**C4 GW_R GND 4.29F
**C3 NET289 GND 1.1F
**C2 NET083 GND 0.5F
**C1 NET088 GND 1.1F
**C0 NET141 GND 0.7F
**C54 NET90 GND 0.45F
**C18 WLPCD0 GND 4F
.ENDS S1100W8_IO_RWCTRL_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IORWBLK_M8                                                           *
* LAST TIME SAVED: DEC 14 17:21:00 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IORWBLK_M8 BLEQB Q DL DLB AWTI BIST BWEB BWEBM D DCLK DM GW_RB WLP
XDIN AWTD BWEB_M NET42 BIST BWEB BWEBM D DM S1100W8_DIN
XSA Q AWTD AWTI DL DLB PGB PREB SAE S1100W8_SA
XIO_WRIN DL DLB NET42 DCLK_DATA NET041 WPG S1100W8_IO_WRIN_M8
XIO_RWCTRL BLEQB NET041 DCLK_DATA PGB PREB SAE WPG BWEB_M DCLK GW_RB WLP
+S1100W8_IO_RWCTRL_M8
**C3 WPG GND 1.7F
**C2 SAE GND 3F
**C8 NET041 GND 1.5F
**C4 PGB GND 4.3F
**C0 DCLK_DATA GND 4.7F
**C5 PREB GND 2.1F
**C7 AWTD GND 1.7F
**C6 BWEB_M GND 1.7F
**C1 NET42 GND 1.7F
.ENDS S1100W8_IORWBLK_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IOYPASS_M8                                                           *
* LAST TIME SAVED: DEC 14 17:22:46 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IOYPASS_M8 BL BLB DL DLB BLEQB YSEL
**C19 NET47 GND 0.97F
*MN0 BL YSEL DL GND NCH W=0.8U L=0.06U
MN0 BL YSEL DL GND NCH W=0.89U L=0.06U
*MN1 BLB YSEL DLB GND NCH W=0.8U L=0.06U
MN1 BLB YSEL DLB GND NCH W=0.89U L=0.06U
MP2 BLB BLEQB BL VDD PCH W=2U L=0.06U
MP0 BL NET47 DL VDD PCH W=0.8U L=0.06U
MP3 VDD BLEQB BLB VDD PCH W=2U L=0.06U
MP1 BLB NET47 DLB VDD PCH W=0.8U L=0.06U
MP4 BL BLEQB VDD VDD PCH W=2U L=0.06U
XI9 NET47 YSEL S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.24U
.ENDS S1100W8_IOYPASS_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_M8                                                                *
* LAST TIME SAVED: DEC  2 19:25:13 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IO_M8 Q BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] BLB[1]
+BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] AWTI BIST_BUF BWEB BWEBM D DCLK DM
+GW_RB WLP Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0]
**CI6_7 YSEL[7] GND 1.7F
**CI6_6 YSEL[6] GND 1.7F
**CI6_5 YSEL[5] GND 1.7F
**CI6_4 YSEL[4] GND 1.7F
**CI6_3 YSEL[3] GND 1.7F
**CI6_2 YSEL[2] GND 1.7F
**CI6_1 YSEL[1] GND 1.7F
**CI6_0 YSEL[0] GND 1.7F
**CI7 NET31 GND 13F
**CI9 NET32 GND 8.13F
**CI11 NET33 GND 8.09F
XI2 NET31 Q NET33 NET32 AWTI BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP S1100W8_IORWBLK_M8
XYSELX4_1 YSEL[7] YSEL[6] YSEL[5] YSEL[4] Y10[3] Y10[2] Y10[1] Y10[0] Y32[1]
+S1100W8_YSELX4
XYSELX4_0 YSEL[3] YSEL[2] YSEL[1] YSEL[0] Y10[3] Y10[2] Y10[1] Y10[0] Y32[0]
+S1100W8_YSELX4
XIYPASS_7 BL[7] BLB[7] NET33 NET32 NET31 YSEL[7] S1100W8_IOYPASS_M8
XIYPASS_6 BL[6] BLB[6] NET33 NET32 NET31 YSEL[6] S1100W8_IOYPASS_M8
XIYPASS_5 BL[5] BLB[5] NET33 NET32 NET31 YSEL[5] S1100W8_IOYPASS_M8
XIYPASS_4 BL[4] BLB[4] NET33 NET32 NET31 YSEL[4] S1100W8_IOYPASS_M8
XIYPASS_3 BL[3] BLB[3] NET33 NET32 NET31 YSEL[3] S1100W8_IOYPASS_M8
XIYPASS_2 BL[2] BLB[2] NET33 NET32 NET31 YSEL[2] S1100W8_IOYPASS_M8
XIYPASS_1 BL[1] BLB[1] NET33 NET32 NET31 YSEL[1] S1100W8_IOYPASS_M8
XIYPASS_0 BL[0] BLB[0] NET33 NET32 NET31 YSEL[0] S1100W8_IOYPASS_M8
.ENDS S1100W8_IO_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_WRIN_M4                                                           *
* LAST TIME SAVED: DEC 14 16:50:06 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IO_WRIN_M4 DL DLB D DCLK DLEQB WPG
XLH_DCLK_M8 D1B DCLK D S1100W8_LH_DCLK
MP7 DL DLEQB VDD VDD PCH W=1U L=0.07U
MP8 VDD DLEQB DLB VDD PCH W=1U L=0.07U
MN2 VDD D1 D2B VDD PCH W=2.5U L=0.07U
MN0 VDD D1B D2 VDD PCH W=2.5U L=0.07U
MN5 DLB WPG D2B GND NCH W=2.5U L=0.07U
MN4 D2 WPG DL GND NCH W=2.5U L=0.07U
MN3 D2B D1 GND GND NCH W=5U L=0.07U
MN1 D2 D1B GND GND NCH W=5U L=0.07U
XI69 D1 D1B S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
**C11 D1B GND 5.983F
**C6 D1 GND 3.851F
**C7 D2B GND 2.669F
**C8 D2 GND 3.188F
.ENDS S1100W8_IO_WRIN_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_RWCTRL_M4                                                         *
* LAST TIME SAVED: DEC 14 16:50:07 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IO_RWCTRL_M4 BLEQB DLEQB DLH PGB PREB SAE WPG BWEB DCLK GW_RB WLP
X_LH_BWEB BWEB_SU DLH BWEB S1100W8_LH_BWEB
XI289 PREB NET0100 NET161 S1100W8_SNOR LP1=0.07U WP1=1.2U LP2=0.07U WP2=1.2U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI288 NET161 WLPCD2 NET163 S1100W8_SNOR LP1=0.07U WP1=0.35U LP2=0.07U WP2=0.35U LN2=0.07U
+WN2=0.3U LN1=0.07U WN1=0.3U
XI249 WPG GW_R NET089 S1100W8_SNOR LP1=0.07U WP1=1.0U LP2=0.07U WP2=1.0U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI133 NET073 WLPCD0 NET_110 GW_R S1100W8_SNAND3 LP3=0.07U WP3=1.75U LP2=0.07U WP2=1.75U
+LP1=0.07U WP1=1.75U LN1=0.07U WN1=1.2U LN2=0.07U WN2=1.2U LN3=0.07U WN3=1.2U
XI250 PGB NET166 GW_R S1100W8_SNAND LP2=0.07U WP2=0.84U LP1=0.07U WP1=0.84U LN1=0.07U
+WN1=0.7U LN2=0.07U WN2=0.7U
XI305 NET90 NET073 WLPCD2 S1100W8_SNAND LP2=0.07U WP2=0.42U LP1=0.07U WP1=0.42U LN1=0.07U
+WN1=0.21U LN2=0.07U WN2=0.21U
XI307 BLEQB WLPCD0 WLPCD4 S1100W8_SNAND LP2=0.07U WP2=1.75U LP1=0.07U WP1=3.5U LN1=0.07U
+WN1=1U LN2=0.07U WN2=1U
XI306 NET289 WLPCD1 BWEB_SU S1100W8_SNAND LP2=0.07U WP2=0.3U LP1=0.07U WP1=0.3U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI339 NET0219 DCLK WLPCD3 S1100W8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI186 NET163 NET93 NET073 S1100W8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI312 NET083 WLPCD0 S1100W8_SINV LP=0.10U WP=0.35U LN=0.10U WN=0.15U
XI73 GW_R GW_RB S1100W8_SINV LP=0.07U WP=1.4U LN=0.07U WN=0.7U
XI348 NET0100 GW_R S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI329 NET0153 WLPCD3 S1100W8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.15U
XI217 WLPCD1 WLPCD0 S1100W8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.28U
XI340 DLH NET0219 S1100W8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.7U
XI287 NET93 NET135 S1100W8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI327 NET141 NET139 S1100W8_SINV LP=0.18U WP=0.35U LN=0.18U WN=0.15U
XI286 NET135 PGB S1100W8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI134 SAE NET073 S1100W8_SINV LP=0.15U WP=0.7U LN=0.1U WN=0.35U
XI321 NET062 NET289 S1100W8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI264 WLPCD4 NET0153 S1100W8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI322 NET089 NET062 S1100W8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.2U
XI185 NET166 NET90 S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.28U
XI299 WLPCD2 NET100 S1100W8_SINV LP=0.07U WP=0.9U LN=0.07U WN=0.3U
XI298 NET100 WLPCD1 S1100W8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI207 NET_110 NET141 S1100W8_SINV LP=0.10U WP=0.7U LN=0.10U WN=0.28U
XI334 DLEQB NET095 S1100W8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
XI337 WLPCD3 WLPCD2 S1100W8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.25U
XI128 WLPCD0 NET085 S1100W8_SINV LP=0.07U WP=1.6U LN=0.07U WN=0.8U
XI315 NET085 WLP S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI333 NET095 BLEQB S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI311 NET088 NET083 S1100W8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
XI310 NET139 NET088 S1100W8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
**C50 WLPCD4 GND 1.317F
**C51 NET135 GND 0.555F
**C17 WLPCD1 GND 1.524F
**C33 NET139 GND 0.850F
**C15 NET0100 GND 2.197F
**C31 NET_110 GND 2.187F
**C13 NET073 GND 3.990F
**C10 NET095 GND 0.690F
**C11 NET0219 GND 1.025F
**C48 WLPCD2 GND 3.190F
**C47 NET166 GND 0.853F
**C26 BWEB_SU GND 2.568F
**C42 NET161 GND 0.935F
**C27 NET93 GND 0.533F
**C43 NET163 GND 1.781F
**C24 NET062 GND 0.737F
**C9 NET0153 GND 1.066F
**C8 WLPCD3 GND 3.831F
**C7 NET100 GND 0.733F
**C6 NET085 GND 1.719F
**C5 NET089 GND 0.959F
**C4 GW_R GND 6.770F
**C3 NET289 GND 0.760F
**C2 NET083 GND 0.902F
**C1 NET088 GND 0.616F
**C0 NET141 GND 0.837F
**C54 NET90 GND 2.157F
**C18 WLPCD0 GND 7.540F
.ENDS S1100W8_IO_RWCTRL_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IORWBLK_M4                                                           *
* LAST TIME SAVED: DEC  8 17:33:56 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IORWBLK_M4 BLEQB Q DL DLB AWTI BIST BWEB BWEBM D DCLK DM GW_RB WLP
XDIN AWTD BWEB_M NET47 BIST BWEB BWEBM D DM S1100W8_DIN
XIO_WRIN DL DLB NET47 DCLK_DATA NET041 WPG S1100W8_IO_WRIN_M4
XIO_RWCTRL BLEQB NET041 DCLK_DATA PGB PREB SAE WPG BWEB_M DCLK GW_RB WLP
+S1100W8_IO_RWCTRL_M4
XSA Q AWTD AWTI DL DLB PGB PREB SAE S1100W8_SA
**C3 WPG GND 3.447F
**C2 SAE GND 5.928F
**C9 BLEQB GND 4.8F
**C8 NET041 GND 1.500F
**C4 PGB GND 6.882F
**C0 DCLK_DATA GND 6.355F
**C5 PREB GND 5.536F
**C6 BWEB_M GND 1.497F
**C7 AWTD GND 6.791F
**C1 NET47 GND 5.644F
.ENDS S1100W8_IORWBLK_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IOYPASS_M4                                                           *
* LAST TIME SAVED: DEC 14 16:50:08 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IOYPASS_M4 BL BLB DL DLB BLEQB YSEL
**C1 NET47 GND 1.979F
*MN0 BL YSEL DL GND NCH W=0.8U L=0.06U
MN0 BL YSEL DL GND NCH W=0.89U L=0.06U
*MN1 BLB YSEL DLB GND NCH W=0.8U L=0.06U
MN1 BLB YSEL DLB GND NCH W=0.89U L=0.06U
MP2 BLB BLEQB BL VDD PCH W=2U L=0.06U
MP0 BL NET47 DL VDD PCH W=0.8U L=0.06U
MP3 VDD BLEQB BLB VDD PCH W=2U L=0.06U
MP1 BLB NET47 DLB VDD PCH W=0.8U L=0.06U
MP4 BL BLEQB VDD VDD PCH W=2U L=0.06U
XI9 NET47 YSEL S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.24U
.ENDS S1100W8_IOYPASS_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_M4                                                                *
* LAST TIME SAVED: DEC 15 14:54:17 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_IO_M4 Q BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] AWTI
+BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP Y10[3] Y10[2] Y10[1] Y10[0]
XI2 NET23 Q NET25 NET24 AWTI BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP S1100W8_IORWBLK_M4
XIYPASS_3 BL[3] BLB[3] NET25 NET24 NET23 Y10[3] S1100W8_IOYPASS_M4
XIYPASS_2 BL[2] BLB[2] NET25 NET24 NET23 Y10[2] S1100W8_IOYPASS_M4
XIYPASS_1 BL[1] BLB[1] NET25 NET24 NET23 Y10[1] S1100W8_IOYPASS_M4
XIYPASS_0 BL[0] BLB[0] NET25 NET24 NET23 Y10[0] S1100W8_IOYPASS_M4
**C4 NET23 GND 15.052F
**C1 NET25 GND 9.518F
**C0 NET24 GND 9.433F
.ENDS S1100W8_IO_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SINV_HVT                                                             *
* LAST TIME SAVED: SEP 21 15:49:08 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_SINV_HVT Y A LP=0.06U WP=0.3U LN=0.06U WN=0.15U
M0 Y A GND GND NCH_HVT W=WN L=LN
M1 VDD A Y VDD PCH_HVT W=WP L=LP
.ENDS S1100W8_SINV_HVT


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V3                                                             *
* LAST TIME SAVED: DEC 14 16:49:42 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_DELAY_V3 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET28 TSEL IN S1100W8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI163 OUT_B NET28 S1100W8_SINV_HVT LP=0.32U WP=0.6U LN=0.32U WN=0.3U
**C153 NET28 GND 0.7F
.ENDS S1100W8_DELAY_V3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V2                                                             *
* LAST TIME SAVED: DEC 14 16:49:31 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_DELAY_V2 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET44 TSEL IN S1100W8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI165 OUT_B NET44 S1100W8_SINV_HVT LP=0.18U WP=0.6U LN=0.18U WN=0.3U
**C153 NET44 GND 0.7F
.ENDS S1100W8_DELAY_V2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V1                                                             *
* LAST TIME SAVED: DEC 14 16:49:18 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_DELAY_V1 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET27 TSEL IN S1100W8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI141 OUT_B NET27 S1100W8_SINV_HVT LP=0.12U WP=0.6U LN=0.12U WN=0.3U
**C151 NET27 GND 1.1F
.ENDS S1100W8_DELAY_V1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_CEB                                                               *
* LAST TIME SAVED: DEC 14 16:50:09 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_LH_CEB Q CP D
XI26 D P2 CP INCP S1100W8_TRANSGATE LP=0.07U WP=1U LN=0.07U WN=1U
MN12 GND Q NET39 GND NCH W=0.15U L=0.07U
MN11 NET39 INCP P2 GND NCH W=0.15U L=0.07U
MP4 NET69 Q VDD VDD PCH W=0.28U L=0.07U
MP5 P2 CP NET69 VDD PCH W=0.28U L=0.07U
XI33 Q P2 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI29 INCP CP S1100W8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
**C1 P2 GND 1.955F
**C0 INCP GND 0.828F
.ENDS S1100W8_LH_CEB


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: PREBUF                                                               *
* LAST TIME SAVED: DEC 14 16:50:09 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_PREBUF SCLK_X SCLK_Y CEB CLK WLPX
X_LH_CEB H1 CK2 NET0309 S1100W8_LH_CEB
XI345 CK2 NET0179 H1 H0 S1100W8_TRANSGATE LP=0.06U WP=3.5U LN=0.06U WN=3.5U
MP4 NET0179 H1 VDD VDD PCH W=2U L=0.06U
XI358 CK2 NET0130 CLK S1100W8_SNOR LP1=0.06U WP1=3U LP2=0.06U WP2=3U LN2=0.06U WN2=3U
+LN1=0.06U WN1=3U
XI356 SCLK_Y NET0179 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=5U M=1
XI382 SCLK_X NET0179 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=5U M=2
XI353 H0 H1 S1100W8_SINV LP=0.06U WP=1U LN=0.06U WN=0.5U
XI354 NET0309 NET0297 S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI357 NET0302 NET0304 S1100W8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI359 NET0304 WLPX S1100W8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI361 NET0130 NET0302 S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI404 NET0297 CEB S1100W8_SINV LP=0.10U WP=0.3U LN=0.10U WN=0.15U
**C8 NET0179 GND 15.756F
**C9 H1 GND 5.364F
**C10 NET0309 GND 1.493F
**C12 H0 GND 1.999F
**C14 NET0297 GND 0.677F
**C39 NET0130 GND 2.062F
**C37 NET0304 GND 0.598F
**C38 NET0302 GND 0.748F
**C43 CK2 GND 7.480F
.ENDS S1100W8_PREBUF


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DFFQ_WEB                                                             *
* LAST TIME SAVED: DEC 14 16:50:10 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_DFFQ_WEB Q CP D
XI30 INV2 P2 INCP CP S1100W8_TRANSGATE LP=0.07U WP=2U LN=0.07U WN=1U
MN17 NET38 Q GND GND NCH W=0.3U L=0.07U
MN15 NET44 INV2 GND GND NCH W=0.2U L=0.07U
MN16 P2 CP NET38 GND NCH W=0.3U L=0.07U
MN14 INV1 INCP NET44 GND NCH W=0.2U L=0.07U
MN13 NET54 D GND GND NCH W=0.3U L=0.07U
MN7 INV1 CP NET54 GND NCH W=0.3U L=0.07U
MP10 NET68 INCP P2 VDD PCH W=0.6U L=0.07U
MP0 VDD D NET78 VDD PCH W=0.6U L=0.07U
MP7 VDD INV2 NET74 VDD PCH W=0.4U L=0.07U
MP6 NET78 INCP INV1 VDD PCH W=0.6U L=0.07U
MP8 NET74 CP INV1 VDD PCH W=0.4U L=0.07U
MP9 VDD Q NET68 VDD PCH W=0.6U L=0.07U
XI31 Q P2 S1100W8_SINV LP=0.07U WP=10U LN=0.07U WN=5U
XI33 INCP CP S1100W8_SINV LP=0.07U WP=1.00U LN=0.07U WN=0.35U
XI29 INV2 INV1 S1100W8_SINV LP=0.07U WP=3.0U LN=0.07U WN=1.5U
**C0 INV1 GND 2.338F
**C1 INCP GND 2.995F
**C2 INV2 GND 2.715F
**C3 P2 GND 5.625F
.ENDS S1100W8_DFFQ_WEB


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CLKBUF                                                               *
* LAST TIME MODIFIED: JULY 24 09:50:10 2006                                       *
*******************************************************************************
.SUBCKT S1100W8_CLKBUF DCLK GW_RB CEB CLK WEB
X_LH_DCLK H3 CK_WEB NET111 S1100W8_LH_DCLK
X_DFFQ_WEB NET69 CK_WEB SH S1100W8_DFFQ_WEB
***------------REMOVE------------------------------------------------------****
**XI273 CLK NET94 H3 H2 TRANSGATE LP=0.06U WP=2.1U LN=0.06U WN=2.1U
**MN10 NET94 H2 GND GND NCH W=0.2U L=0.1U
***------------ADD BELOW MOS------------------------------------------------------****
MP10 DCLK0 H3 VDD VDD PCH W=0.4U L=0.06U
XI1274 NET94 DCLK0 S1100W8_SINV LP=0.06U WP=4U LN=0.06U WN=2U 
MP1 VDD CLK NET001 VDD PCH W=1U L=0.06U
MP2 NET001 H2 DCLK0 VDD PCH W=1U L=0.06U
MN1 NET002 H3 DCLK0 GND NCH W=1U L=0.06U
MN2 GND CLK NET002 GND NCH W=1U L=0.06U
***-----------------------------------------------------------------------------*********
XI271 SH CEB WEB S1100W8_SNOR LP1=0.07U WP1=0.45U LP2=0.07U WP2=0.45U LN2=0.07U WN2=0.15U
+LN1=0.07U WN1=0.15U
XI246 GW_RB NET69 S1100W8_SINV LP=0.06U WP=9U LN=0.06U WN=4.5U M=2
XI280 H2 H3 S1100W8_SINV LP=0.06U WP=0.35U LN=0.06U WN=0.15U
XI277 NET111 SH S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI202 CK_WEB CLK S1100W8_SINV LP=0.06U WP=0.8U LN=0.06U WN=0.8U
XI274 DCLK NET94 S1100W8_SINV LP=0.06U WP=8U LN=0.06U WN=8U M=2
**C43 SH GND 4.641F
**C18 CK_WEB GND 7.391F
**C19 NET69 GND 12.723F
**C21 NET94 GND 13.840F
**C24 H3 GND 4.176F
**C26 NET111 GND 1.130F
**C27 SH GND 4.641F
**C25 H2 GND 1.913F
.ENDS S1100W8_CLKBUF


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M16V1                                                         *
* LAST TIME SAVED: DEC  1 14:30:39 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_WLPGEN_M16V1 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK
+TM TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 NET122 D02 SEL[3] SELN[3] SELN[2] S1100W8_DELAY_V3
XI337 D02 NET122 D01 SEL[2] SELN[2] SELN[1] S1100W8_DELAY_V2
XI326 D01 NET122 NET0214 SEL[1] SELN[1] SELN[0] S1100W8_DELAY_V1
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S1100W8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S1100W8_CLKBUF
**XI324 NET122 NET0214 SEL[0] SELN[0] TRANSGATE LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI324 NET122 NET1227 SEL[0] SELN[0] S1100W8_TRANSGATE LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI238 D1 T0 NET132 CLK_K S1100W8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S1100W8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET169 CLK_KB CLK S1100W8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN7 NET96 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET097 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET096 GND NCH W=5U L=0.06U
MN0 NET096 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET96 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET0198 NET097 GND NCH W=5U L=0.07U
MP5 VDD TME NET0108 VDD PCH W=10U L=0.06U M=2
MP9 NET80 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET0119 NET0198 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET0108 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET80 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET0119 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI219 NET169 WLP_RESET WLPSTART S1100W8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI482 WLP_RESET NET122 NET210 S1100W8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U LN1=0.06U
+WN1=1.0U LN2=0.06U WN2=1.0U
XI328 SELN[0] SEL0N SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S1100W8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI383 NET0198 WLPTEST S1100W8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI386 TRWLPB TRWLP S1100W8_SINV LP=0.2U WP=1.0U LN=0.2U WN=0.4U
XI471 SEL[3] SELN[3] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET0323 S1100W8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET0321 CEB S1100W8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET0348 WLPSTART S1100W8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET0354 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET0354 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI371 NET0323 NET0321 S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI292 NET0214 TRWLPB S1100W8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI283 CLK_KB CLK S1100W8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
**XI493 NET209 NET122 SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI493 NET1227 NET0214 S1100W8_SINV LP=0.06U WP=0.755U LN=0.06U WN=0.2U
XI495 NET213 NET208 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI296 CLK_K NET132 S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI297 NET132 CLK S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**XI494 NET208 NET209 SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI494 NET208 NET122 S1100W8_SINV LP=0.06U WP=0.755U LN=0.06U WN=0.2U
XI473 SEL1 SEL1N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI497 NET210 TRWLP S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI315 TME TMEB S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI496 NET211 NET213 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
**CI414 D03 GND 0.7F
**C36 TRWLPB GND 5.4F
**CI428 D02 GND 1.2F
**C40 NET0354 GND 5.6F
**CI410 SEL0 GND 2.1F
**CI446 TME GND 5.5F
**CI426 D01 GND 1.3F
**CI420 SEL0N GND 2.9F
**CI434 NET0214 GND 1.5F
**CI448 TMEB GND 6.1F
**C0 T2 GND 6.1F
**C4 NET132 GND 0.7F
**CI418 SEL1 GND 2.7F
**C34 WLPSTART GND 13.1F
**C35 NET0348 GND 8.2F
**CI432 NET0198 GND 5.2F
**C30 NET0323 GND 0.7F
**C15 NET0321 GND 0.7F
**CI422 SEL1N GND 2.8F
**C32 D1 GND 1.4F
**C1 T1 GND 3.2F
**C5 CLK_K GND 0.8F
**CI444 SELN[0] GND 3.9F
**C22 CLK_KB GND 2.2F
**CI442 SEL[0] GND 4.1F
**C33 T0 GND 1.0F
**C31 NET169 GND 5.6F
**C2 WLP_RESET GND 5.5F
.ENDS S1100W8_WLPGEN_M16V1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CEBBISMX                                                             *
* LAST TIME SAVED: NOV 30 14:35:28 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_CEBBISMX MXOUT A AM BISTC BISTT
**C0 GND NET30 1.033F
XI5 MXOUT NET30 S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
MP15 Z21 BISTT NET30 VDD PCH W=0.5U L=0.06U
MP14 VDD A Z21 VDD PCH W=0.5U L=0.06U
MP7 VDD AM Z22 VDD PCH W=0.5U L=0.06U
MP6 Z22 BISTC NET30 VDD PCH W=0.5U L=0.06U
MN15 NET30 BISTC Z23 GND NCH W=0.25U L=0.06U
MN14 NET30 BISTT Z24 GND NCH W=0.25U L=0.06U
MN13 Z23 A GND GND NCH W=0.25U L=0.06U
MN6 Z24 AM GND GND NCH W=0.25U L=0.06U
.ENDS S1100W8_CEBBISMX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AWTD_M16                                                             *
* LAST TIME SAVED: OCT  4 16:21:02 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_AWTD_M16 AWTI AWT
XINV0 AWTI Z1 S1100W8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI9 Z1 AWT S1100W8_SINV LP=0.07U WP=3U LN=0.07U WN=1.5U
.ENDS S1100W8_AWTD_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISTD_M16                                                            *
* LAST TIME SAVED: OCT  4 16:22:00 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BISTD_M16 BISTC BISTT BIST
XI13 BISTT BISTC S1100W8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI14 BISTC BIST S1100W8_SINV LP=0.07U WP=3.2U LN=0.07U WN=1.6U
.ENDS S1100W8_BISTD_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISIN_M16                                                            *
* LAST TIME SAVED: DEC  1 14:16:28 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BISIN_M16 AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM
XCEBMX CEBX CEB CEBM BISTC BIST_BUF S1100W8_CEBBISMX
XWEBMX WEBX WEB WEBM BISTC BIST_BUF S1100W8_CEBBISMX
XAWTD AWTI AWT S1100W8_AWTD_M16
XBISTD BISTC BIST_BUF BIST S1100W8_BISTD_M16
.ENDS S1100W8_BISIN_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SRAM_TIEL                                                            *
* LAST TIME SAVED: MAY 16 14:03:38 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_SRAM_TIEL Z
XI49 Z NET14 S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=4U
MN1 GND NET14 NET32 GND NCH W=0.15U L=0.07U
MN0 NET32 NET32 GND GND NCH W=0.15U L=0.07U
MP0 VDD NET32 NET14 VDD PCH W=0.3U L=0.07U
.ENDS S1100W8_SRAM_TIEL


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_YPD_M16                                                           *
* LAST TIME SAVED: SEP 30 15:10:52 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_LH_YPD_M16 Q CP D
XI26 D P2 INCPN CP S1100W8_TRANSGATE LP=0.07U WP=2U LN=0.07U WN=2U
MN0 GND Q NET38 GND NCH W=0.2U L=0.07U
MN1 NET38 CP P2 GND NCH W=0.2U L=0.07U
MP4 NET49 Q VDD VDD PCH W=0.5U L=0.07U
MP5 P2 INCPN NET49 VDD PCH W=0.5U L=0.07U
XI23 Q P2 S1100W8_SINV LP=0.07U WP=8U LN=0.07U WN=4U
XI29 INCPN CP S1100W8_SINV LP=0.07U WP=1.2U LN=0.07U WN=0.6U
**C2 P2 GND 3F
**C3 INCPN GND 1.5F
.ENDS S1100W8_LH_YPD_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPRE10_M16                                                           *
* LAST TIME SAVED: DEC 13 14:07:14 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_YPRE10_M16 Y10[3] Y10[2] Y10[1] Y10[0] BISTT SCLK Y[1] Y[0] YM[1] YM[0]
MP0 NET43 BISTC Y1N VDD PCH W=0.3U L=0.07U
MP15 NET40 BISTT Y0N VDD PCH W=0.3U L=0.07U
MP14 VDD Y[0] NET40 VDD PCH W=0.3U L=0.07U
MP7 VDD YM[0] NET31 VDD PCH W=0.3U L=0.07U
MP6 NET31 BISTC Y0N VDD PCH W=0.3U L=0.07U
MP1 VDD YM[1] NET43 VDD PCH W=0.3U L=0.07U
MP2 VDD Y[1] NET22 VDD PCH W=0.3U L=0.07U
MP3 NET22 BISTT Y1N VDD PCH W=0.3U L=0.07U
MN3 Y1N BISTC NET46 GND NCH W=0.15U L=0.07U
MN2 Y1N BISTT NET49 GND NCH W=0.15U L=0.07U
MN15 Y0N BISTC NET55 GND NCH W=0.15U L=0.07U
MN14 Y0N BISTT NET52 GND NCH W=0.15U L=0.07U
MN13 NET55 Y[0] GND GND NCH W=0.15U L=0.07U
MN6 NET52 YM[0] GND GND NCH W=0.15U L=0.07U
MN0 NET49 YM[1] GND GND NCH W=0.15U L=0.07U
MN1 NET46 Y[1] GND GND NCH W=0.15U L=0.07U
XLH_YPD_3 Y10[3] SCLK NET073 S1100W8_LH_YPD_M16
XLH_YPD_2 Y10[2] SCLK NET075 S1100W8_LH_YPD_M16
XLH_YPD_0 Y10[0] SCLK NET070 S1100W8_LH_YPD_M16
XLH_YPD_1 Y10[1] SCLK NET083 S1100W8_LH_YPD_M16
XI154 NET35 Y0N DY[1] S1100W8_SNAND LP2=0.06U WP2=0.18U LP1=0.06U WP1=0.18U LN1=0.06U
+WN1=0.2U LN2=0.06U WN2=0.2U
XI152 NET036 DY[0] Y1N S1100W8_SNAND LP2=0.06U WP2=0.18U LP1=0.06U WP1=0.18U LN1=0.06U
+WN1=0.2U LN2=0.06U WN2=0.2U
XI39 NET41 Y0N Y1N S1100W8_SNAND LP2=0.06U WP2=0.18U LP1=0.06U WP1=0.18U LN1=0.06U WN1=0.2U
+LN2=0.06U WN2=0.2U
XI153 NET53 DY[0] DY[1] S1100W8_SNAND LP2=0.06U WP2=0.18U LP1=0.06U WP1=0.18U LN1=0.06U
+WN1=0.2U LN2=0.06U WN2=0.2U
XI5 DY[0] Y0N S1100W8_SINV LP=0.07U LN=0.07U
XI579 DY[1] Y1N S1100W8_SINV LP=0.07U LN=0.07U
XI200 NET073 NET077 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI199 NET075 NET088 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI123 NET072 NET41 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI124 NET070 NET072 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI202 NET088 NET35 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI190 NET083 NET090 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI201 NET090 NET036 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI215 BISTC BISTT S1100W8_SINV LP=0.07U LN=0.07U
XI203 NET077 NET53 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
**C36 Y1N GND 2F
**C28 DY[0] GND 1.3F
**C27 DY[1] GND 1.3F
**C29 Y0N GND 2F
**C13 NET35 GND 0.5F
**C14 NET088 GND 0.5F
**C15 NET077 GND 0.5F
**C12 NET53 GND 0.5F
**C16 NET090 GND 0.5F
**C17 NET072 GND 0.5F
**C10 NET41 GND 0.5F
**C18 NET070 GND 0.5F
**C19 NET083 GND 0.5F
**C20 NET073 GND 0.5F
**C21 NET075 GND 0.5F
**C11 NET036 GND 0.5F
.ENDS S1100W8_YPRE10_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPREDEC_M16                                                          *
* LAST TIME SAVED: SEP 30 16:22:48 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_YPREDEC_M16 Y10[3] Y10[2] Y10[1] Y10[0] BISTT SCLK Y[1] Y[0] YM[1]
+YM[0]
XYPRE10 Y10[3] Y10[2] Y10[1] Y10[0] BISTT SCLK Y[1] Y[0] YM[1] YM[0] S1100W8_YPRE10_M16
.ENDS S1100W8_YPREDEC_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_XPD8                                                              *
* LAST TIME SAVED: DEC 14 17:25:05 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_LH_XPD8 Q CP D
XI26 NET043 P1 INCPN CP S1100W8_TRANSGATE LP=0.07U WP=3U LN=0.07U WN=1.5U
MN12 GND Q NET39 GND NCH W=0.25U L=0.07U
MN11 NET39 NET042 P1 GND NCH W=0.25U L=0.07U
MP4 NET69 Q VDD VDD PCH W=0.5U L=0.07U
MP5 P1 INCPN NET69 VDD PCH W=0.5U L=0.07U
XI38 NET042 INCPN S1100W8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.15U
XI24 Q P1 S1100W8_SINV LP=0.07U WP=6U LN=0.07U WN=3U M=2
XI29 INCPN CP S1100W8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.5U
XI36 NET043 D S1100W8_SINV LP=0.07U WP=3U LN=0.07U WN=1.5U
**C1 INCPN GND 2.759F
**C0 P1 GND 10.654F
**C39 NET042 GND 0.780F
**C3 NET043 GND 3.343F
.ENDS S1100W8_LH_XPD8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XPRE8                                                                *
* LAST TIME SAVED: DEC 14 17:24:55 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_XPRE8 XPRE[7] XPRE[6] XPRE[5] XPRE[4] XPRE[3] XPRE[2] XPRE[1] XPRE[0]
+BIST WLP X[2] X[1] X[0] XM[2] XM[1] XM[0]
MP9 NET51 BISTC X2N VDD PCH W=0.5U L=0.06U
MP0 NET48 BISTC X1N VDD PCH W=0.5U L=0.06U
MP1 VDD X[1] NET39 VDD PCH W=0.5U L=0.06U
MP2 VDD XM[1] NET48 VDD PCH W=0.5U L=0.06U
MP3 NET39 BISTT X1N VDD PCH W=0.5U L=0.06U
MP6 NET36 BISTT X0N VDD PCH W=0.5U L=0.06U
MP7 VDD XM[0] NET27 VDD PCH W=0.5U L=0.06U
MP10 VDD X[0] NET36 VDD PCH W=0.5U L=0.06U
MP11 NET27 BISTC X0N VDD PCH W=0.5U L=0.06U
MP5 VDD X[2] NET60 VDD PCH W=0.5U L=0.06U
MP8 VDD XM[2] NET51 VDD PCH W=0.5U L=0.06U
MP4 NET60 BISTT X2N VDD PCH W=0.5U L=0.06U
MN0 NET84 X[1] GND GND NCH W=0.25U L=0.06U
MN1 NET81 XM[1] GND GND NCH W=0.25U L=0.06U
MN2 X1N BISTC NET84 GND NCH W=0.25U L=0.06U
MN3 X1N BISTT NET81 GND NCH W=0.25U L=0.06U
MN7 NET87 X[2] GND GND NCH W=0.25U L=0.06U
MN8 NET90 XM[2] GND GND NCH W=0.25U L=0.06U
MN4 X2N BISTC NET87 GND NCH W=0.25U L=0.06U
MN6 X0N BISTT NET66 GND NCH W=0.25U L=0.06U
MN9 X0N BISTC NET63 GND NCH W=0.25U L=0.06U
MN10 NET66 XM[0] GND GND NCH W=0.25U L=0.06U
MN11 NET63 X[0] GND GND NCH W=0.25U L=0.06U
MN5 X2N BISTT NET90 GND NCH W=0.25U L=0.06U
XLH_XPD8_2 XPRE[2] WLP NET162 S1100W8_LH_XPD8
XLH_XPD8_3 XPRE[3] WLP NET097 S1100W8_LH_XPD8
XLH_XPD8_7 XPRE[7] WLP NET085 S1100W8_LH_XPD8
XLH_XPD8_5 XPRE[5] WLP NET156 S1100W8_LH_XPD8
XLH_XPD8_1 XPRE[1] WLP NET165 S1100W8_LH_XPD8
XLH_XPD8_6 XPRE[6] WLP NET171 S1100W8_LH_XPD8
XLH_XPD8_0 XPRE[0] WLP NET089 S1100W8_LH_XPD8
XLH_XPD8_4 XPRE[4] WLP NET153 S1100W8_LH_XPD8
XI624 BISTT BISTC S1100W8_SINV LP=0.06U LN=0.06U
XI582 NET165 NET038 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI608 X1 X1N S1100W8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI447 NET089 NET167 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI590 NET156 NET046 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI584 NET097 NET050 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI588 X2 X2N S1100W8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI615 X0 X0N S1100W8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI591 NET171 NET026 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI592 NET085 NET034 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI583 NET162 NET054 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI589 NET153 NET030 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI623 BISTC BIST S1100W8_SINV LP=0.06U LN=0.06U
XI600 NET030 X0N X1N X2 S1100W8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI602 NET026 X0N X1 X2 S1100W8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI598 NET054 X0N X1 X2N S1100W8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI603 NET034 X0 X1 X2 S1100W8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI599 NET050 X0 X1 X2N S1100W8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI597 NET038 X0 X1N X2N S1100W8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI407 NET167 X0N X1N X2N S1100W8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI601 NET046 X0 X1N X2 S1100W8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
**C71 BISTT GND 4.975F
**C72 BISTC GND 5.774F
**C57 NET046 GND 1.321F
**C58 NET030 GND 1.363F
**C67 X1 GND 3.655F
**C68 X1N GND 4.286F
**C66 X2N GND 4.779F
**C46 NET038 GND 1.346F
**C63 NET085 GND 3.233F
**C64 NET156 GND 3.230F
**C65 NET153 GND 3.332F
**C47 NET054 GND 1.329F
**C59 NET165 GND 3.192F
**C50 NET050 GND 1.314F
**C32 X2 GND 3.573F
**C69 X0N GND 6.023F
**C70 X0 GND 5.270F
**C40 NET089 GND 3.244F
**C44 NET167 GND 1.348F
**C60 NET097 GND 3.231F
**C61 NET162 GND 3.239F
**C62 NET171 GND 3.306F
**C55 NET034 GND 1.349F
**C56 NET026 GND 1.307F
.ENDS S1100W8_XPRE8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XPREDEC888                                                           *
* LAST TIME SAVED: DEC  5 14:42:50 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_XPREDEC888 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1]
+XPD0[0] XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0]
+XPD2[7] XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLK
+X[8] X[7] X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4]
+XM[3] XM[2] XM[1] XM[0]
XPRE8_A XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+BIST_BUF SCLK X[2] X[1] X[0] XM[2] XM[1] XM[0] S1100W8_XPRE8
XPRE8_B XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0]
+BIST_BUF SCLK X[5] X[4] X[3] XM[5] XM[4] XM[3] S1100W8_XPRE8
XPRE8_C XPD2[7] XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0]
+BIST_BUF SCLK X[8] X[7] X[6] XM[8] XM[7] XM[6] S1100W8_XPRE8
.ENDS S1100W8_XPREDEC888


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL888_M16                                                          *
* LAST TIME SAVED: DEC  1 14:30:43 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_CTRL888_M16 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7]
+XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2] Y10[1]
+Y10[0] Y32[3] Y32[2] Y32[1] Y32[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1]
+TSEL[0] WEB WEBM WLPTEST X[8] X[7] X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[8]
+XM[7] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0] Y[3] Y[2] Y[1] Y[0] YM[3]
+YM[2] YM[1] YM[0]
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S1100W8_WLPGEN_M16V1
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S1100W8_BISIN_M16
XI180 CTRL_TIEL S1100W8_SRAM_TIEL
XI182 CTRL_TIELB S1100W8_SRAM_TIEL
XYPREDEC32 Y32[3] Y32[2] Y32[1] Y32[0] BIST_BUF NET65 Y[3] Y[2] YM[3] YM[2]
+S1100W8_YPREDEC_M16
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S1100W8_YPREDEC_M16
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[7]
+XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7] XPD2[6]
+XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[8] X[7] X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1]
+XM[0] S1100W8_XPREDEC888
.ENDS S1100W8_CTRL888_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M8V1                                                          *
* LAST TIME SAVED: DEC 14 17:41:43 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_WLPGEN_M8V1 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK TM
+TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 PRE_WLP_RESET D02 SEL[3] SELN[3] SELN[2] S1100W8_DELAY_V3
XI337 D02 PRE_WLP_RESET D01 SEL[2] SELN[2] SELN[1] S1100W8_DELAY_V2
XI326 D01 PRE_WLP_RESET TRWLPBB SEL[1] SELN[1] SELN[0] S1100W8_DELAY_V1
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S1100W8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S1100W8_CLKBUF
XI238 D1 T0 NET259 CLK_K S1100W8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S1100W8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET148 CLK_KB CLK S1100W8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN4 NET151 TRWLPBB GND GND NCH W=0.5U L=0.06U
MN5 PRE_WLP_RESET SEL[0] NET151 GND NCH W=0.5U L=0.06U
MN7 NET165 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET155 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET161 GND NCH W=5U L=0.06U
MN0 NET161 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET165 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET227 NET155 GND NCH W=5U L=0.07U
MP7 NET175 SELN[0] PRE_WLP_RESET VDD PCH W=1.0U L=0.06U
MP10 VDD TRWLPBB NET175 VDD PCH W=1.0U L=0.06U M=1
MP5 VDD TME NET179 VDD PCH W=10U L=0.06U M=2
MP9 NET173 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET186 NET227 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET179 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET173 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET186 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI482 WLP_RESET PRE_WLP_RESET NET217 S1100W8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U
+LN1=0.06U WN1=1.0U LN2=0.06U WN2=1.0U
XI219 NET148 WLP_RESET WLPSTART S1100W8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI328 SELN[0] SEL0N SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S1100W8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI477 NET227 WLPTEST S1100W8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI495 NET209 NET210 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI507 TRWLPBB TRWLPB S1100W8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI494 NET210 NET215 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI386 TRWLPB TRWLP S1100W8_SINV LP=0.12U WP=1.0U LN=0.12U WN=0.4U
XI496 NET218 NET209 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI493 NET215 PRE_WLP_RESET S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI471 SEL[3] SELN[3] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET253 S1100W8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET251 CEB S1100W8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET239 WLPSTART S1100W8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET239 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET243 NET239 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET243 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET239 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI371 NET253 NET251 S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI497 NET217 TRWLP S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI283 CLK_KB CLK S1100W8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
XI296 CLK_K NET259 S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI297 NET259 CLK S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI473 SEL1 SEL1N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI315 TME TMEB S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**C47 SELN[0] GND 2.7F
**C48 SEL[0] GND 2.7F
**C49 SELN[2] GND 2.7F
**C50 SEL[2] GND 2.7F
**C44 SEL[3] GND 2.7F
**C36 TRWLPB GND 5.4F
**C428 D02 GND 1.2F
**C40 NET243 GND 5.6F
**C410 SEL0 GND 2.1F
**C446 TME GND 5.5F
**C426 D01 GND 1.3F
**C420 SEL0N GND 2.9F
**C448 TMEB GND 6.1F
**C0 T2 GND 6.1F
**C4 NET259 GND 0.7F
**C418 SEL1 GND 2.7F
**C34 WLPSTART GND 13.1F
**C35 NET239 GND 8.2F
**C432 NET227 GND 5.2F
**C30 NET253 GND 0.7F
**C43 SELN[3] GND 2.7F
**C29 NET251 GND 0.6F
**C422 SEL1N GND 2.8F
**C32 D1 GND 1.4F
**C1 T1 GND 3.2F
**C5 CLK_K GND 0.8F
**C2 WLP_RESET GND 5.5F
**C430 PRE_WLP_RESET GND 4.2F
**C45 SELN[1] GND 2.7F
**C22 CLK_KB GND 2.2F
**C33 T0 GND 1.0F
**C46 SEL[1] GND 2.7F
**C31 NET148 GND 5.6F
**C51 TRWLPBB GND 5.4F
.ENDS S1100W8_WLPGEN_M8V1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AWTD_M8                                                              *
* LAST TIME SAVED: OCT  4 10:09:37 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_AWTD_M8 AWTI AWT
XINV0 AWTI Z1 S1100W8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI9 Z1 AWT S1100W8_SINV LP=0.07U WP=3U LN=0.07U WN=1.5U
.ENDS S1100W8_AWTD_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISTD_M8                                                             *
* LAST TIME SAVED: OCT  4 10:38:52 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BISTD_M8 BISTC BISTT BIST
XI13 BISTT BISTC S1100W8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI14 BISTC BIST S1100W8_SINV LP=0.07U WP=3.2U LN=0.07U WN=1.6U
.ENDS S1100W8_BISTD_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISIN_M8                                                             *
* LAST TIME SAVED: DEC  1 14:10:29 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BISIN_M8 AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM
XCEBMX CEBX CEB CEBM BISTC BIST_BUF S1100W8_CEBBISMX
XWEBMX WEBX WEB WEBM BISTC BIST_BUF S1100W8_CEBBISMX
XAWTD AWTI AWT S1100W8_AWTD_M8
XBISTD BISTC BIST_BUF BIST S1100W8_BISTD_M8
.ENDS S1100W8_BISIN_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_YPD_M8                                                            *
* LAST TIME SAVED: MAY 25 14:13:06 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_LH_YPD_M8 Q CP D
XI26 D P2 INCPN CP S1100W8_TRANSGATE LP=0.07U WP=2U LN=0.07U WN=2U
MN0 GND Q NET38 GND NCH W=0.2U L=0.07U
MN1 NET38 CP P2 GND NCH W=0.2U L=0.07U
MP4 NET49 Q VDD VDD PCH W=0.5U L=0.07U
MP5 P2 INCPN NET49 VDD PCH W=0.5U L=0.07U
XI23 Q P2 S1100W8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI29 INCPN CP S1100W8_SINV LP=0.07U WP=1.2U LN=0.07U WN=0.6U
**C2 P2 GND 3.9F
**C3 INCPN GND 1.5F
.ENDS S1100W8_LH_YPD_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPRE10_M2                                                            *
* LAST TIME SAVED: SEP 29 14:55:40 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_YPRE10_M2 Y32[1] Y32[0] BISTT SCLK Y[0] YM[0]
MP14 VDD Y[0] Z21 VDD PCH W=0.3U L=0.07U
MP15 Z21 BISTT Y0N VDD PCH W=0.3U L=0.07U
MP7 VDD YM[0] Z22 VDD PCH W=0.3U L=0.07U
MP6 Z22 BISTC Y0N VDD PCH W=0.3U L=0.07U
MN15 Y0N BISTC Z23 GND NCH W=0.15U L=0.07U
MN14 Y0N BISTT Z24 GND NCH W=0.15U L=0.07U
MN6 Z24 YM[0] GND GND NCH W=0.15U L=0.07U
MN13 Z23 Y[0] GND GND NCH W=0.15U L=0.07U
XLH_YPD_0 Y32[0] SCLK NET070 S1100W8_LH_YPD_M8
XLH_YPD_1 Y32[1] SCLK NET083 S1100W8_LH_YPD_M8
XI5 Y0 Y0N S1100W8_SINV LP=0.07U LN=0.07U
XI123 NET072 NET41 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI124 NET070 NET072 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI201 NET083 NET090 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI205 BISTC BISTT S1100W8_SINV LP=0.07U LN=0.07U
XI199 NET41 Y0N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI202 NET090 NET036 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI203 NET036 Y0 S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
**C28 Y0 GND 0.7F
**C29 Y0N GND 1.1F
**C16 NET090 GND 1.1F
**C17 NET072 GND 1.1F
**C10 NET41 GND 1.6F
**C18 NET070 GND 2.9F
**C19 NET083 GND 2.9F
**C11 NET036 GND 1.6F
.ENDS S1100W8_YPRE10_M2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPREDEC_M2                                                           *
* LAST TIME SAVED: OCT 24 09:46:40 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_YPREDEC_M2 Y32[1] Y32[0] BIST_BUF SCLK Y[0] YM[0]
XYPRE10 Y32[1] Y32[0] BIST_BUF SCLK Y[0] YM[0] S1100W8_YPRE10_M2
.ENDS S1100W8_YPREDEC_M2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPRE10_M8                                                            *
* LAST TIME SAVED: OCT  4 10:00:07 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_YPRE10_M8 Y10[3] Y10[2] Y10[1] Y10[0] BISTT SCLK Y[1] Y[0] YM[1] YM[0]
MN3 Y1N BISTC NET44 GND NCH W=0.15U L=0.07U
MN2 Y1N BISTT NET173 GND NCH W=0.15U L=0.07U
MN15 Y0N BISTC NET174 GND NCH W=0.15U L=0.07U
MN14 Y0N BISTT NET38 GND NCH W=0.15U L=0.07U
MN13 NET174 Y[0] GND GND NCH W=0.15U L=0.07U
MN6 NET38 YM[0] GND GND NCH W=0.15U L=0.07U
MN0 NET173 YM[1] GND GND NCH W=0.15U L=0.07U
MN1 NET44 Y[1] GND GND NCH W=0.15U L=0.07U
MP0 NET47 BISTC Y1N VDD PCH W=0.3U L=0.07U
MP15 NET50 BISTT Y0N VDD PCH W=0.3U L=0.07U
MP14 VDD Y[0] NET50 VDD PCH W=0.3U L=0.07U
MP7 VDD YM[0] NET59 VDD PCH W=0.3U L=0.07U
MP6 NET59 BISTC Y0N VDD PCH W=0.3U L=0.07U
MP1 VDD YM[1] NET47 VDD PCH W=0.3U L=0.07U
MP2 VDD Y[1] NET68 VDD PCH W=0.3U L=0.07U
MP3 NET68 BISTT Y1N VDD PCH W=0.3U L=0.07U
XLH_YPD_3 Y10[3] SCLK NET073 S1100W8_LH_YPD_M8
XLH_YPD_2 Y10[2] SCLK NET075 S1100W8_LH_YPD_M8
XLH_YPD_0 Y10[0] SCLK NET070 S1100W8_LH_YPD_M8
XLH_YPD_1 Y10[1] SCLK NET083 S1100W8_LH_YPD_M8
XI211 NET35 Y0N DY[1] S1100W8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI210 NET036 DY[0] Y1N S1100W8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI212 NET53 DY[0] DY[1] S1100W8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI39 NET41 Y0N Y1N S1100W8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI215 BISTC BISTT S1100W8_SINV LP=0.07U LN=0.07U
XI5 DY[0] Y0N S1100W8_SINV LP=0.07U LN=0.07U
XI579 DY[1] Y1N S1100W8_SINV LP=0.07U LN=0.07U
XI202 NET075 NET088 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI201 NET083 NET090 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI123 NET072 NET41 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI124 NET070 NET072 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI206 NET077 NET53 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI203 NET073 NET077 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI205 NET088 NET35 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI204 NET090 NET036 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
**C36 Y1N GND 2F
**C28 DY[0] GND 1.3F
**C27 DY[1] GND 1.3F
**C29 Y0N GND 2F
**C13 NET35 GND 1.3F
**C14 NET088 GND 1.1F
**C15 NET077 GND 1.1F
**C12 NET53 GND 1.3F
**C16 NET090 GND 1.1F
**C17 NET072 GND 1.1F
**C10 NET41 GND 1.3F
**C18 NET070 GND 2.8F
**C19 NET083 GND 2.8F
**C20 NET073 GND 2.8F
**C21 NET075 GND 2.8F
**C11 NET036 GND 1.3F
.ENDS S1100W8_YPRE10_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPREDEC_M8                                                           *
* LAST TIME SAVED: OCT 24 09:46:40 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_YPREDEC_M8 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF SCLK Y[1] Y[0] YM[1]
+YM[0]
XYPRE10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF SCLK Y[1] Y[0] YM[1] YM[0]
+S1100W8_YPRE10_M8
.ENDS S1100W8_YPREDEC_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL888_M8                                                           *
* LAST TIME SAVED: DEC 14 17:41:45 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_CTRL888_M8 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7]
+XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2] Y10[1]
+Y10[0] Y32[1] Y32[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1] TSEL[0] WEB WEBM
+WLPTEST X[8] X[7] X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5]
+XM[4] XM[3] XM[2] XM[1] XM[0] Y[2] Y[1] Y[0] YM[2] YM[1] YM[0]
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S1100W8_WLPGEN_M8V1
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S1100W8_BISIN_M8
XSRM_TIEL CTRL_TIEL S1100W8_SRAM_TIEL
XSRM_TIEL2 CTRL_TIELB S1100W8_SRAM_TIEL
**C184 SCLKX GND 34.2F
**C187 NET65 GND 15.3F
**C7 WEBX GND 3.022F
XYPREDEC32 Y32[1] Y32[0] BIST_BUF NET65 Y[2] YM[2] S1100W8_YPREDEC_M2
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S1100W8_YPREDEC_M8
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[7]
+XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7] XPD2[6]
+XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[8] X[7] X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1]
+XM[0] S1100W8_XPREDEC888
.ENDS S1100W8_CTRL888_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M4V1                                                          *
* LAST TIME SAVED: DEC 14 16:49:46 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_WLPGEN_M4V1 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK TM
+TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 NET170 D02 SEL[3] SELN[3] SELN[2] S1100W8_DELAY_V3
XI337 D02 NET170 D01 SEL[2] SELN[2] SELN[1] S1100W8_DELAY_V2
XI326 D01 NET170 NET0214 SEL[1] SELN[1] SELN[0] S1100W8_DELAY_V1
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S1100W8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S1100W8_CLKBUF
XI238 D1 T0 NET132 CLK_K S1100W8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S1100W8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET169 CLK_KB CLK S1100W8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN4 NET333 NET0214 GND GND NCH W=0.5U L=0.06U
MN5 NET170 SEL[0] NET333 GND NCH W=0.5U L=0.06U
MN7 NET96 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET097 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET096 GND NCH W=5U L=0.06U
MN0 NET096 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET96 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET0198 NET097 GND NCH W=5U L=0.07U
MP10 VDD NET0214 NET173 VDD PCH W=1.0U L=0.06U M=1
MP5 VDD TME NET0108 VDD PCH W=10U L=0.06U M=2
MP7 NET173 SELN[0] NET170 VDD PCH W=1.0U L=0.06U
MP9 NET80 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET0119 NET0198 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET0108 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET80 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET0119 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI219 NET169 WLP_RESET WLPSTART S1100W8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI482 WLP_RESET NET170 NET218 S1100W8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U LN1=0.06U
+WN1=1.0U LN2=0.06U WN2=1.0U
XI328 SELN[0] SEL0N SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S1100W8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI383 NET0198 WLPTEST S1100W8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI386 TRWLPB TRWLP S1100W8_SINV LP=0.12U WP=1.0U LN=0.12U WN=0.4U
XI496 NET219 NET226 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI494 NET224 NET220 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI471 SEL[3] SELN[3] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET0323 S1100W8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET0321 CEB S1100W8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET0348 WLPSTART S1100W8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET0354 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET0354 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI493 NET220 NET170 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI371 NET0323 NET0321 S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI292 NET0214 TRWLPB S1100W8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI283 CLK_KB CLK S1100W8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
XI296 CLK_K NET132 S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI497 NET218 TRWLP S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI495 NET226 NET224 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI297 NET132 CLK S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI473 SEL1 SEL1N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI315 TME TMEB S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**C36 TRWLPB GND 3.009F
**C44 NET170 GND 5.266F
**C428 D02 GND 1.950F
**C40 NET0354 GND 13.839F
**C43 WLP_RESET GND 4.630F
**C410 SEL0 GND 2.687F
**C446 TME GND 11.753F
**C426 D01 GND 2.319F
**C420 SEL0N GND 2.317F
**C434 NET0214 GND 3.637F
**C448 TMEB GND 11.368F
**C0 T2 GND 9.532F
**C4 NET132 GND 1.008F
**C418 SEL1 GND 2.583F
**C34 WLPSTART GND 28.916F
**C35 NET0348 GND 25.077F
**C432 NET0198 GND 6.135F
**C30 NET0323 GND 1.326F
**C29 NET0321 GND 0.782F
**C422 SEL1N GND 2.592F
**C32 D1 GND 1.821F
**C1 T1 GND 5.899F
**C5 CLK_K GND 1.749F
**C22 CLK_KB GND 6.158F
**C33 T0 GND 3.232F
**C31 NET169 GND 2.156F
.ENDS S1100W8_WLPGEN_M4V1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AWTD_M4                                                              *
* LAST TIME SAVED: DEC 14 16:50:10 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_AWTD_M4 AWTI AWT
**C0 Z1 GND 8.034F
XINV0 AWTI Z1 S1100W8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI9 Z1 AWT S1100W8_SINV LP=0.07U WP=3U LN=0.07U WN=1.5U
.ENDS S1100W8_AWTD_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISTD_M4                                                             *
* LAST TIME SAVED: OCT 13 22:07:21 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BISTD_M4 BISTC BIST_BUF BIST
XI13 BIST_BUF BISTC S1100W8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI14 BISTC BIST S1100W8_SINV LP=0.07U WP=3.2U LN=0.07U WN=1.6U
.ENDS S1100W8_BISTD_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISIN_M4                                                             *
* LAST TIME SAVED: DEC 14 19:54:47 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BISIN_M4 AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM
XCEBMX CEBX CEB CEBM BISTC BIST_BUF S1100W8_CEBBISMX
XWEBMX WEBX WEB WEBM BISTC BIST_BUF S1100W8_CEBBISMX
**C0 BISTC GND 9.597F
XAWTD AWTI AWT S1100W8_AWTD_M4
XBISTD BISTC BIST_BUF BIST S1100W8_BISTD_M4
.ENDS S1100W8_BISIN_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_YPD_M4                                                            *
* LAST TIME SAVED: NOV 10 11:38:58 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_LH_YPD_M4 Q CP D
XI26 D P2 INCPN CP S1100W8_TRANSGATE LP=0.07U WP=2U LN=0.07U WN=2U
MN0 GND Q NET38 GND NCH W=0.2U L=0.07U
MN1 NET38 CP P2 GND NCH W=0.2U L=0.07U
MP4 NET49 Q VDD VDD PCH W=0.5U L=0.07U
MP5 P2 INCPN NET49 VDD PCH W=0.5U L=0.07U
XI23 Q P2 S1100W8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI29 INCPN CP S1100W8_SINV LP=0.07U WP=1.2U LN=0.07U WN=0.6U
**C2 P2 GND 13.447F
**C3 INCPN GND 2.178F
.ENDS S1100W8_LH_YPD_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPRE10_M4                                                            *
* LAST TIME SAVED: DEC 14 16:50:11 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_YPRE10_M4 Y10[3] Y10[2] Y10[1] Y10[0] BIST SCLK Y[1] Y[0] YM[1] YM[0]
XLH_YPD_3 Y10[3] SCLK NET073 S1100W8_LH_YPD_M4
XLH_YPD_2 Y10[2] SCLK NET075 S1100W8_LH_YPD_M4
XLH_YPD_0 Y10[0] SCLK NET070 S1100W8_LH_YPD_M4
XLH_YPD_1 Y10[1] SCLK NET083 S1100W8_LH_YPD_M4
MN3 Y1N BISTC NET44 GND NCH W=0.15U L=0.07U
MN2 Y1N BISTT NET173 GND NCH W=0.15U L=0.07U
MN15 Y0N BISTC NET174 GND NCH W=0.15U L=0.07U
MN14 Y0N BISTT NET38 GND NCH W=0.15U L=0.07U
MN13 NET174 Y[0] GND GND NCH W=0.15U L=0.07U
MN6 NET38 YM[0] GND GND NCH W=0.15U L=0.07U
MN0 NET173 YM[1] GND GND NCH W=0.15U L=0.07U
MN1 NET44 Y[1] GND GND NCH W=0.15U L=0.07U
MP0 NET47 BISTC Y1N VDD PCH W=0.3U L=0.07U
MP15 NET50 BISTT Y0N VDD PCH W=0.3U L=0.07U
MP14 VDD Y[0] NET50 VDD PCH W=0.3U L=0.07U
MP7 VDD YM[0] NET59 VDD PCH W=0.3U L=0.07U
MP6 NET59 BISTC Y0N VDD PCH W=0.3U L=0.07U
MP1 VDD YM[1] NET47 VDD PCH W=0.3U L=0.07U
MP2 VDD Y[1] NET68 VDD PCH W=0.3U L=0.07U
MP3 NET68 BISTT Y1N VDD PCH W=0.3U L=0.07U
XI211 NET35 Y0N DY[1] S1100W8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI210 NET036 DY[0] Y1N S1100W8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI212 NET53 DY[0] DY[1] S1100W8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI39 NET41 Y0N Y1N S1100W8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI217 BISTT BISTC S1100W8_SINV LP=0.07U LN=0.07U
XI215 BISTC BIST S1100W8_SINV LP=0.07U LN=0.07U
XI5 DY[0] Y0N S1100W8_SINV LP=0.07U LN=0.07U
XI579 DY[1] Y1N S1100W8_SINV LP=0.07U LN=0.07U
XI202 NET075 NET088 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI201 NET083 NET090 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI123 NET072 NET41 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI124 NET070 NET072 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI206 NET077 NET53 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI203 NET073 NET077 S1100W8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI205 NET088 NET35 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI204 NET090 NET036 S1100W8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
**C26 BISTC GND 3.305F
**C30 BISTT GND 2.787F
**C36 Y1N GND 3.008F
**C28 DY[0] GND 1.800F
**C27 DY[1] GND 1.800F
**C29 Y0N GND 3.177F
**C13 NET35 GND 1.134F
**C14 NET088 GND 1.642F
**C15 NET077 GND 1.516F
**C12 NET53 GND 1.460F
**C16 NET090 GND 1.796F
**C17 NET072 GND 1.425F
**C10 NET41 GND 1.330F
**C18 NET070 GND 2.637F
**C19 NET083 GND 2.970F
**C20 NET073 GND 2.854F
**C21 NET075 GND 2.503F
**C11 NET036 GND 1.426F
.ENDS S1100W8_YPRE10_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPREDEC_M4                                                           *
* LAST TIME SAVED: OCT 13 22:07:22 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_YPREDEC_M4 Y10[3] Y10[2] Y10[1] Y10[0] BIST SCLK Y[1] Y[0] YM[1] YM[0]
XYPRE10 Y10[3] Y10[2] Y10[1] Y10[0] BIST SCLK Y[1] Y[0] YM[1] YM[0] S1100W8_YPRE10_M4
.ENDS S1100W8_YPREDEC_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL888_M4                                                           *
* LAST TIME SAVED: DEC 14 17:10:45 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_CTRL888_M4 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7]
+XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2] Y10[1]
+Y10[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1] TSEL[0] WEB WEBM WLPTEST X[8]
+X[7] X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4] XM[3]
+XM[2] XM[1] XM[0] Y[1] Y[0] YM[1] YM[0]
**C5 NET241 GND 12.589F
**C6 SCLKX GND 58.558F
**C7 WEBX GND 3.022F
XCTRL_WLPGEN DCLK GW_RB SCLKX NET241 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S1100W8_WLPGEN_M4V1
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S1100W8_BISIN_M4
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET241 Y[1] Y[0] YM[1] YM[0]
+S1100W8_YPREDEC_M4
XI180 CTRL_TIEL S1100W8_SRAM_TIEL
XI182 CTRL_TIELB S1100W8_SRAM_TIEL
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[7]
+XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7] XPD2[6]
+XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[8] X[7] X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1]
+XM[0] S1100W8_XPREDEC888
.ENDS S1100W8_CTRL888_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V6                                                             *
* LAST TIME SAVED: DEC 14 15:09:57 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_DELAY_V6 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET28 TSEL IN S1100W8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI163 OUT_B NET28 S1100W8_SINV_HVT LP=0.16U WP=0.6U LN=0.16U WN=0.3U
**CI153 NET28 GND 0.7F
.ENDS S1100W8_DELAY_V6


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V5                                                             *
* LAST TIME SAVED: DEC 14 15:09:45 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_DELAY_V5 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET44 TSEL IN S1100W8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI165 OUT_B NET44 S1100W8_SINV_HVT LP=0.06U WP=0.6U LN=0.06U WN=0.3U
**CI153 NET44 GND 0.7F
.ENDS S1100W8_DELAY_V5


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V4                                                             *
* LAST TIME SAVED: DEC 15 14:54:17 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_DELAY_V4 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET27 TSEL IN S1100W8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI141 OUT_B NET27 S1100W8_SINV_HVT LP=0.06U WP=0.6U LN=0.06U WN=0.3U
**C151 NET27 GND 0.946F
.ENDS S1100W8_DELAY_V4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M16V3                                                         *
* LAST TIME SAVED: DEC  1 14:40:33 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_WLPGEN_M16V3 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK
+TM TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 NET122 D02 SEL[3] SELN[3] SELN[2] S1100W8_DELAY_V6
XI337 D02 NET122 D01 SEL[2] SELN[2] SELN[1] S1100W8_DELAY_V5
XI326 D01 NET122 NET0214 SEL[1] SELN[1] SELN[0] S1100W8_DELAY_V4
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S1100W8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S1100W8_CLKBUF
**XI324 NET122 NET0214 SEL[0] SELN[0] TRANSGATE LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI324 NET122 NET1227 SEL[0] SELN[0] S1100W8_TRANSGATE LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI238 D1 T0 NET132 CLK_K S1100W8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S1100W8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET169 CLK_KB CLK S1100W8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN7 NET96 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET097 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET096 GND NCH W=5U L=0.06U
MN0 NET096 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET96 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET0198 NET097 GND NCH W=5U L=0.07U
MP5 VDD TME NET0108 VDD PCH W=10U L=0.06U M=2
MP9 NET80 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET0119 NET0198 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET0108 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET80 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET0119 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI219 NET169 WLP_RESET WLPSTART S1100W8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI482 WLP_RESET NET122 NET210 S1100W8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U LN1=0.06U
+WN1=1.0U LN2=0.06U WN2=1.0U
XI328 SELN[0] SEL0N SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S1100W8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI383 NET0198 WLPTEST S1100W8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI386 TRWLPB TRWLP S1100W8_SINV LP=0.2U WP=1.0U LN=0.2U WN=0.4U
XI471 SEL[3] SELN[3] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET0323 S1100W8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET0321 CEB S1100W8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET0348 WLPSTART S1100W8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET0354 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET0354 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI371 NET0323 NET0321 S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI292 NET0214 TRWLPB S1100W8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI283 CLK_KB CLK S1100W8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
**XI493 NET209 NET122 SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI493 NET1227 NET0214 S1100W8_SINV LP=0.06U WP=0.755U LN=0.06U WN=0.2U
XI495 NET213 NET208 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI296 CLK_K NET132 S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI297 NET132 CLK S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**XI494 NET208 NET209 SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI494 NET208 NET122 S1100W8_SINV LP=0.06U WP=0.755U LN=0.06U WN=0.2U
XI473 SEL1 SEL1N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI497 NET210 TRWLP S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI315 TME TMEB S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI496 NET211 NET213 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
**CI414 D03 GND 0.7F
**C36 TRWLPB GND 5.4F
**CI428 D02 GND 1.2F
**C40 NET0354 GND 5.6F
**CI410 SEL0 GND 2.1F
**CI446 TME GND 5.5F
**CI426 D01 GND 1.3F
**CI420 SEL0N GND 2.9F
**CI434 NET0214 GND 1.5F
**CI448 TMEB GND 6.1F
**C0 T2 GND 6.1F
**C4 NET132 GND 0.7F
**CI418 SEL1 GND 2.7F
**C34 WLPSTART GND 13.1F
**C35 NET0348 GND 8.2F
**CI432 NET0198 GND 5.2F
**C30 NET0323 GND 0.7F
**C29 NET0321 GND 0.6F
**CI422 SEL1N GND 2.8F
**C32 D1 GND 1.4F
**C1 T1 GND 3.2F
**C5 CLK_K GND 0.8F
**CI444 SELN[0] GND 3.9F
**C22 CLK_KB GND 2.2F
**CI442 SEL[0] GND 4.1F
**C33 T0 GND 1.0F
**C31 NET169 GND 5.6F
**C2 WLP_RESET GND 5.5F
.ENDS S1100W8_WLPGEN_M16V3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XPRE4                                                                *
* LAST TIME SAVED: DEC 14 15:46:20 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_XPRE4 XPRE[3] XPRE[2] XPRE[1] XPRE[0] BIST WLP X[1] X[0] XM[1] XM[0]
MN11 NET41 X[0] GND GND NCH W=0.25U L=0.06U
MN10 NET38 XM[0] GND GND NCH W=0.25U L=0.06U
MN9 X0N BISTC NET41 GND NCH W=0.25U L=0.06U
MN6 X0N BISTT NET38 GND NCH W=0.25U L=0.06U
MN3 X1N BISTT NET23 GND NCH W=0.25U L=0.06U
MN2 X1N BISTC NET20 GND NCH W=0.25U L=0.06U
MN1 NET23 XM[1] GND GND NCH W=0.25U L=0.06U
MN0 NET20 X[1] GND GND NCH W=0.25U L=0.06U
MP11 NET65 BISTC X0N VDD PCH W=0.5U L=0.06U
MP10 VDD X[0] NET56 VDD PCH W=0.5U L=0.06U
MP7 VDD XM[0] NET65 VDD PCH W=0.5U L=0.06U
MP6 NET56 BISTT X0N VDD PCH W=0.5U L=0.06U
MP3 NET53 BISTT X1N VDD PCH W=0.5U L=0.06U
MP2 VDD XM[1] NET44 VDD PCH W=0.5U L=0.06U
MP1 VDD X[1] NET53 VDD PCH W=0.5U L=0.06U
MP0 NET44 BISTC X1N VDD PCH W=0.5U L=0.06U
XLH_XPD8_2 XPRE[2] WLP NET162 S1100W8_LH_XPD8
XLH_XPD8_3 XPRE[3] WLP NET097 S1100W8_LH_XPD8
XLH_XPD8_1 XPRE[1] WLP NET165 S1100W8_LH_XPD8
XLH_XPD8_0 XPRE[0] WLP NET089 S1100W8_LH_XPD8
XI582 BISTT BISTC S1100W8_SINV LP=0.06U LN=0.06U
XI575 NET165 NET038 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.31U
XI623 BISTC BIST S1100W8_SINV LP=0.06U LN=0.06U
XI615 X0 X0N S1100W8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI608 X1 X1N S1100W8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI447 NET089 NET167 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.31U
XI577 NET097 NET050 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.31U
XI576 NET162 NET054 S1100W8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.31U
XI574 NET050 X0 X1 S1100W8_SNAND LP2=0.07U WP2=0.15U LP1=0.07U WP1=0.15U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI572 NET038 X0 X1N S1100W8_SNAND LP2=0.07U WP2=0.15U LP1=0.07U WP1=0.15U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI573 NET054 X0N X1 S1100W8_SNAND LP2=0.07U WP2=0.15U LP1=0.07U WP1=0.15U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI407 NET167 X0N X1N S1100W8_SNAND LP2=0.07U WP2=0.15U LP1=0.07U WP1=0.15U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
**C70 X0 GND 1.483F
**C69 X0N GND 3.380F
**C68 X1N GND 2.374F
**C67 X1 GND 1.667F
**C46 NET038 GND 1.453F
**C47 NET054 GND 1.481F
**C59 NET165 GND 3.147F
**C50 NET050 GND 1.384F
**C40 NET089 GND 3.277F
**C44 NET167 GND 1.470F
**C60 NET097 GND 3.216F
**C61 NET162 GND 3.122F
.ENDS S1100W8_XPRE4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XPREDEC844                                                           *
* LAST TIME SAVED: DEC  6 09:48:41 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_XPREDEC844 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1]
+XPD0[0] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST
+SCLK X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1]
+XM[0]
XPRE4_B XPD1[3] XPD1[2] XPD1[1] XPD1[0] BIST SCLK X[4] X[3] XM[4] XM[3] S1100W8_XPRE4
XPRE4_C XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST SCLK X[6] X[5] XM[6] XM[5] S1100W8_XPRE4
XPRE8_A XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] BIST
+SCLK X[2] X[1] X[0] XM[2] XM[1] XM[0] S1100W8_XPRE8
.ENDS S1100W8_XPREDEC844


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL844_M16                                                          *
* LAST TIME SAVED: DEC  1 14:18:20 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_CTRL844_M16 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2]
+Y10[1] Y10[0] Y32[3] Y32[2] Y32[1] Y32[0] AWT BIST CEB CEBM CLK TM TRWLP
+TSEL[1] TSEL[0] WEB WEBM WLPTEST X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[6]
+XM[5] XM[4] XM[3] XM[2] XM[1] XM[0] Y[3] Y[2] Y[1] Y[0] YM[3] YM[2] YM[1]
+YM[0]
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S1100W8_WLPGEN_M16V3
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S1100W8_BISIN_M16
XI180 CTRL_TIEL S1100W8_SRAM_TIEL
XI182 CTRL_TIELB S1100W8_SRAM_TIEL
XYPREDEC32 Y32[3] Y32[2] Y32[1] Y32[0] BIST_BUF NET65 Y[3] Y[2] YM[3] YM[2]
+S1100W8_YPREDEC_M16
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S1100W8_YPREDEC_M16
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[3]
+XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0]
+S1100W8_XPREDEC844
.ENDS S1100W8_CTRL844_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M8V3                                                          *
* LAST TIME SAVED: DEC 14 19:38:34 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_WLPGEN_M8V3 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK TM
+TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 PRE_WLP_RESET D02 SEL[3] SELN[3] SELN[2] S1100W8_DELAY_V6
XI337 D02 PRE_WLP_RESET D01 SEL[2] SELN[2] SELN[1] S1100W8_DELAY_V5
XI326 D01 PRE_WLP_RESET TRWLPBB SEL[1] SELN[1] SELN[0] S1100W8_DELAY_V4
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S1100W8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S1100W8_CLKBUF
XI238 D1 T0 NET259 CLK_K S1100W8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S1100W8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET148 CLK_KB CLK S1100W8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN4 NET151 TRWLPBB GND GND NCH W=0.5U L=0.06U
MN5 PRE_WLP_RESET SEL[0] NET151 GND NCH W=0.5U L=0.06U
MN7 NET165 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET155 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET161 GND NCH W=5U L=0.06U
MN0 NET161 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET165 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET227 NET155 GND NCH W=5U L=0.07U
MP7 NET175 SELN[0] PRE_WLP_RESET VDD PCH W=1.0U L=0.06U
MP10 VDD TRWLPBB NET175 VDD PCH W=1.0U L=0.06U M=1
MP5 VDD TME NET179 VDD PCH W=10U L=0.06U M=2
MP9 NET173 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET186 NET227 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET179 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET173 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET186 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI482 WLP_RESET PRE_WLP_RESET NET217 S1100W8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U
+LN1=0.06U WN1=1.0U LN2=0.06U WN2=1.0U
XI219 NET148 WLP_RESET WLPSTART S1100W8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI328 SELN[0] SEL0N SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S1100W8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI477 NET227 WLPTEST S1100W8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI495 NET209 NET210 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI507 TRWLPBB TRWLPB S1100W8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI494 NET210 NET215 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI386 TRWLPB TRWLP S1100W8_SINV LP=0.12U WP=1.0U LN=0.12U WN=0.4U
XI496 NET218 NET209 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI493 NET215 PRE_WLP_RESET S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI471 SEL[3] SELN[3] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET253 S1100W8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET251 CEB S1100W8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET239 WLPSTART S1100W8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET239 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET243 NET239 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET243 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET239 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI371 NET253 NET251 S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI497 NET217 TRWLP S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI283 CLK_KB CLK S1100W8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
XI296 CLK_K NET259 S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI297 NET259 CLK S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI473 SEL1 SEL1N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI315 TME TMEB S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**C47 SELN[0] GND 2.7F
**C48 SEL[0] GND 2.7F
**C49 SELN[2] GND 2.7F
**C50 SEL[2] GND 2.7F
**C44 SEL[3] GND 2.7F
**C36 TRWLPB GND 5.4F
**CI428 D02 GND 1.2F
**C40 NET243 GND 5.6F
**CI410 SEL0 GND 2.1F
**CI446 TME GND 5.5F
**CI426 D01 GND 1.3F
**CI420 SEL0N GND 2.9F
**CI448 TMEB GND 6.1F
**C0 T2 GND 6.1F
**C4 NET259 GND 0.7F
**CI418 SEL1 GND 2.7F
**C34 WLPSTART GND 13.1F
**C35 NET239 GND 8.2F
**CI432 NET227 GND 5.2F
**C30 NET253 GND 0.7F
**C43 SELN[3] GND 2.7F
**C15 NET251 GND 0.7F
**CI422 SEL1N GND 2.8F
**C32 D1 GND 1.4F
**C1 T1 GND 3.2F
**C5 CLK_K GND 0.8F
**C2 WLP_RESET GND 5.5F
**CI430 PRE_WLP_RESET GND 4.2F
**C45 SELN[1] GND 2.7F
**C22 CLK_KB GND 2.2F
**C33 T0 GND 1.0F
**C46 SEL[1] GND 2.7F
**C31 NET148 GND 5.6F
**C51 TRWLPBB GND 5.4F
.ENDS S1100W8_WLPGEN_M8V3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL844_M8                                                           *
* LAST TIME SAVED: DEC 14 19:38:13 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_CTRL844_M8 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2]
+Y10[1] Y10[0] Y32[1] Y32[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1] TSEL[0] WEB
+WEBM WLPTEST X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2]
+XM[1] XM[0] Y[2] Y[1] Y[0] YM[2] YM[1] YM[0]
**C16 BIST_BUF GND 29.489F
**C5 NET65 GND 12.844F
**C6 SCLKX GND 42.727F
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S1100W8_WLPGEN_M8V3
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S1100W8_BISIN_M8
XI180 CTRL_TIEL S1100W8_SRAM_TIEL
XI182 CTRL_TIELB S1100W8_SRAM_TIEL
XYPREDEC32 Y32[1] Y32[0] BIST_BUF NET65 Y[2] YM[2] S1100W8_YPREDEC_M2
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S1100W8_YPREDEC_M8
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[3]
+XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0]
+S1100W8_XPREDEC844
.ENDS S1100W8_CTRL844_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M4V3                                                          *
* LAST TIME SAVED: DEC 14 16:35:44 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_WLPGEN_M4V3 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK TM
+TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 NET170 D02 SEL[3] SELN[3] SELN[2] S1100W8_DELAY_V6
XI337 D02 NET170 D01 SEL[2] SELN[2] SELN[1] S1100W8_DELAY_V5
XI326 D01 NET170 NET0214 SEL[1] SELN[1] SELN[0] S1100W8_DELAY_V4
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S1100W8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S1100W8_CLKBUF
XI238 D1 T0 NET132 CLK_K S1100W8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S1100W8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET169 CLK_KB CLK S1100W8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN4 NET333 NET0214 GND GND NCH W=0.5U L=0.06U
MN5 NET170 SEL[0] NET333 GND NCH W=0.5U L=0.06U
MN7 NET96 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET097 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET096 GND NCH W=5U L=0.06U
MN0 NET096 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET96 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET0198 NET097 GND NCH W=5U L=0.07U
MP10 VDD NET0214 NET173 VDD PCH W=1.0U L=0.06U M=1
MP5 VDD TME NET0108 VDD PCH W=10U L=0.06U M=2
MP7 NET173 SELN[0] NET170 VDD PCH W=1.0U L=0.06U
MP9 NET80 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET0119 NET0198 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET0108 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET80 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET0119 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI219 NET169 WLP_RESET WLPSTART S1100W8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI482 WLP_RESET NET170 NET218 S1100W8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U LN1=0.06U
+WN1=1.0U LN2=0.06U WN2=1.0U
XI328 SELN[0] SEL0N SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S1100W8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S1100W8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI383 NET0198 WLPTEST S1100W8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI386 TRWLPB TRWLP S1100W8_SINV LP=0.12U WP=1.0U LN=0.12U WN=0.4U
XI496 NET219 NET226 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI494 NET224 NET220 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI471 SEL[3] SELN[3] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET0323 S1100W8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET0321 CEB S1100W8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET0348 WLPSTART S1100W8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET0354 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET0354 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET0348 S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S1100W8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI493 NET220 NET170 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI371 NET0323 NET0321 S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI292 NET0214 TRWLPB S1100W8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI283 CLK_KB CLK S1100W8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
XI296 CLK_K NET132 S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI497 NET218 TRWLP S1100W8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI495 NET226 NET224 S1100W8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI297 NET132 CLK S1100W8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI473 SEL1 SEL1N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S1100W8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI315 TME TMEB S1100W8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**C36 TRWLPB GND 3.301F
**C428 D02 GND 1.848F
**C40 NET0354 GND 13.287F
**C43 WLP_RESET GND 4.827F
**C410 SEL0 GND 2.559F
**C446 TME GND 11.593F
**C426 D01 GND 2.144F
**C420 SEL0N GND 2.663F
**C434 NET0214 GND 3.842F
**C448 TMEB GND 11.386F
**C0 T2 GND 10.101F
**C4 NET132 GND 0.992F
**C418 SEL1 GND 2.410F
**C34 WLPSTART GND 29.449F
**C35 NET0348 GND 25.222F
**CI432 NET0198 GND 5.2F
**C30 NET0323 GND 1.156F
**C15 NET0321 GND 0.780F
**C422 SEL1N GND 2.768F
**C32 D1 GND 1.699F
**C1 T1 GND 5.839F
**C5 CLK_K GND 1.716F
**C22 CLK_KB GND 6.404F
**C33 T0 GND 3.299F
**C31 NET169 GND 2.481F
.ENDS S1100W8_WLPGEN_M4V3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL844_M4                                                           *
* LAST TIME SAVED: DEC 14 15:38:03 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_CTRL844_M4 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2]
+Y10[1] Y10[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1] TSEL[0] WEB WEBM WLPTEST
+X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0]
+Y[1] Y[0] YM[1] YM[0]
**C7 WEBX GND 2.856F
**C16 BIST_BUF GND 29.489F
**C6 SCLKX GND 42.727F
**C5 NET65 GND 12.844F
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S1100W8_WLPGEN_M4V3
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S1100W8_BISIN_M4
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S1100W8_YPREDEC_M4
XI180 CTRL_TIEL S1100W8_SRAM_TIEL
XI182 CTRL_TIELB S1100W8_SRAM_TIEL
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[3]
+XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0]
+S1100W8_XPREDEC844
.ENDS S1100W8_CTRL844_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MDEC_TRK                                                             *
* LAST TIME SAVED: DEC 14 16:50:12 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_MDEC_TRK WLOUT WLPY WLPYB
XI280 WLOUT NET21 S1100W8_SINV_HVTP LN=0.06U WN=5U    LP=0.07U WP=10U    M=2
XI290 NET33 NET15 S1100W8_SINV LP=0.06U WP=0.8U  LN=0.06U WN=0.8U 
MN2 NET15 NET25 GND GND NCH W=0.5U L=0.06U
MN0 NET21 NET33 WLPY GND NCH W=2.0U   L=0.06U
MN1 NET20 NET20 GND GND NCH W=0.5U L=0.06U
MP0 VDD NET33 NET21 VDD PCH W=2.0U   L=0.06U
MP1 NET21 WLPYB VDD VDD PCH W=2.0U      L=0.06U
MP2 VDD NET20 NET25 VDD PCH W=1U L=0.06U
**C3 NET21 GND 9.553F
**C4 NET33 GND 3.064F
.ENDS S1100W8_MDEC_TRK


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BCELL                                                                *
* LAST TIME SAVED: OCT 19 14:40:20 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_BCELL BL BLB WL
MN1 BL_IN BLB_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U  AD=0.02P AS=0.011P PD=0.6U
+PS=0.3U
MN5 GND BL_IN BLB_IN GND NCHPD_HVTSR W=0.14U  L=0.065U  AD=0.02P AS=0.011P PD=0.6U
+PS=0.3U
MN3 BL WL BL_IN GND NCHPG_HVTSR W=0.09U  L=0.075U AD=0.02P AS=0.008P PD=0.6U PS=0.275U
MN0 BLB_IN WL BLB GND NCHPG_HVTSR W=0.09U  L=0.075U AD=0.02P AS=0.008P PD=0.6U
+PS=0.275U
MP2 VDD BL_IN BLB_IN VDD PCHPU_HVTSR W=0.08U  L=0.065U  AD=0.009P AS=0.008P PD=0.34U
+PS=0.265U
MP0 BL_IN BLB_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U  AD=0.009P AS=0.008P PD=0.34U
+PS=0.265U
**C1 BL_IN GND 0.15F
**C0 BLB_IN GND 0.15F
.ENDS S1100W8_BCELL


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CELLX4                                                               *
* LAST TIME SAVED: MAY 17 15:57:24 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_CELLX4 BL[0] BL[1] BLB[0] BLB[1] WL[0] WL[1]
XI7 BLB[1] BL[1] WL[1] S1100W8_BCELL
XBCELL1 BLB[1] BL[1] WL[0] S1100W8_BCELL
XI6 BLB[0] BL[0] WL[1] S1100W8_BCELL
XBCELL0 BLB[0] BL[0] WL[0] S1100W8_BCELL
.ENDS S1100W8_CELLX4


*******************************************************************************
* MAIN CIRCUIT NETLIST:                                                       *
*                                                                             *
* BLOCK: LEAFCELL                                                             *
* LAST TIME SAVED: DEC 15 15:43:07 2005                                       *
*******************************************************************************
.SUBCKT S1100W8_LEAFCELL
XI25 NET183[0] NET183[1] NET184 NET185 NET182[0] NET182[1] S1100W8_TRKDUMX2
XI24 NET187[0] NET187[1] NET189 NET190 NET188 NET186[0] NET186[1] S1100W8_TRKNORX2
XI23 NET192[0] NET192[1] NET101 NET195 NET193 NET191[0] NET191[1] S1100W8_TRKMINX2
XI3 NET11 NET412 NET486 NET8 NET7 S1100W8_TRKMIN
XI4 NET6 NET4 NET459 NET13 NET22 NET23 S1100W8_TRKNOR
XI2 NET17 NET15 NET492 NET442 NET12 S1100W8_TRKDUM
XI21 NET473 S1100W8_SRAM_TIEH
XI17 NET0306[0] NET0306[1] NET0306[2] NET0306[3] NET268 NET315 NET260
+NET0305[0] NET0305[1] NET0305[2] NET0305[3] NET312 NET281 S1100W8_XDRVX2
XI8 NET155 NET147[0] NET147[1] NET147[2] NET147[3] NET147[4] NET147[5]
+NET147[6] NET147[7] NET147[8] NET147[9] NET147[10] NET147[11] NET147[12]
+NET147[13] NET147[14] NET147[15] NET146[0] NET146[1] NET146[2] NET146[3]
+NET146[4] NET146[5] NET146[6] NET146[7] NET146[8] NET146[9] NET146[10]
+NET146[11] NET146[12] NET146[13] NET146[14] NET146[15] NET254 NET330 NET154
+NET252 NET153 NET152 NET253 NET151 NET149 NET148[0] NET148[1] NET148[2]
+NET148[3] NET145[0] NET145[1] NET145[2] NET145[3] S1100W8_IO_M16
XI7 NET166 NET156[0] NET156[1] NET156[2] NET156[3] NET156[4] NET156[5]
+NET156[6] NET156[7] NET157[0] NET157[1] NET157[2] NET157[3] NET157[4]
+NET157[5] NET157[6] NET157[7] NET269 NET221 NET165 NET267 NET164 NET163 NET266
+NET162 NET160 NET159[0] NET159[1] NET159[2] NET159[3] NET158[0] NET158[1]
+S1100W8_IO_M8
XI6 NET174 NET175[0] NET175[1] NET175[2] NET175[3] NET176[0] NET176[1]
+NET176[2] NET176[3] NET280 NET194 NET173 NET282 NET172 NET171 NET45 NET170
+NET168 NET167[0] NET167[1] NET167[2] NET167[3] S1100W8_IO_M4
XI14 NET300 NET334 NET381 NET229 NET216 NET213 NET20 NET19 NET18 NET203
+NET207[0] NET207[1] NET207[2] NET207[3] NET207[4] NET207[5] NET207[6]
+NET207[7] NET325[0] NET325[1] NET325[2] NET325[3] NET325[4] NET325[5]
+NET325[6] NET325[7] NET326[0] NET326[1] NET326[2] NET326[3] NET326[4]
+NET326[5] NET326[6] NET326[7] NET208[0] NET208[1] NET208[2] NET208[3]
+NET214[0] NET214[1] NET214[2] NET214[3] NET296 NET295 NET223 NET299 NET201
+NET224 NET217 NET211[0] NET211[1] NET220 NET294 NET112 NET324[0] NET324[1]
+NET324[2] NET324[3] NET324[4] NET324[5] NET324[6] NET324[7] NET324[8]
+NET293[0] NET293[1] NET293[2] NET293[3] NET293[4] NET293[5] NET293[6]
+NET293[7] NET293[8] NET219[0] NET219[1] NET219[2] NET219[3] NET297[0]
+NET297[1] NET297[2] NET297[3] S1100W8_CTRL888_M16
XI13 NET331 NET144 NET405 NET415 NET72 NET71 NET69 NET68 NET67 NET66 NET65[0]
+NET65[1] NET65[2] NET65[3] NET65[4] NET65[5] NET65[6] NET65[7] NET349[0]
+NET349[1] NET349[2] NET349[3] NET349[4] NET349[5] NET349[6] NET349[7]
+NET350[0] NET350[1] NET350[2] NET350[3] NET350[4] NET350[5] NET350[6]
+NET350[7] NET62[0] NET62[1] NET62[2] NET62[3] NET51[0] NET51[1] NET64 NET70
+NET61 NET328 NET60 NET58 NET57 NET56[0] NET56[1] NET55 NET327 NET233 NET348[0]
+NET348[1] NET348[2] NET348[3] NET348[4] NET348[5] NET348[6] NET348[7]
+NET348[8] NET332[0] NET332[1] NET332[2] NET332[3] NET332[4] NET332[5]
+NET332[6] NET332[7] NET332[8] NET49[0] NET49[1] NET49[2] NET333[0] NET333[1]
+NET333[2] S1100W8_CTRL888_M8
XI12 NET364 NET234 NET431 NET401 NET120 NET119 NET117 NET116 NET115 NET114
+NET113[0] NET113[1] NET113[2] NET113[3] NET113[4] NET113[5] NET113[6]
+NET113[7] NET375[0] NET375[1] NET375[2] NET375[3] NET375[4] NET375[5]
+NET375[6] NET375[7] NET374[0] NET374[1] NET374[2] NET374[3] NET374[4]
+NET374[5] NET374[6] NET374[7] NET110[0] NET110[1] NET110[2] NET110[3] NET362
+NET363 NET109 NET359 NET108 NET106 NET105 NET104[0] NET104[1] NET103 NET357
+NET205 NET373[0] NET373[1] NET373[2] NET373[3] NET373[4] NET373[5] NET373[6]
+NET373[7] NET373[8] NET360[0] NET360[1] NET360[2] NET360[3] NET360[4]
+NET360[5] NET360[6] NET360[7] NET360[8] NET99[0] NET99[1] NET361[0] NET361[1]
+S1100W8_CTRL888_M4
XI11 NET395 NET414 NET455 NET413 NET47 NET46 NET44 NET43 NET42 NET41 NET40[0]
+NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] NET40[6] NET40[7] NET39[0]
+NET39[1] NET39[2] NET39[3] NET38[0] NET38[1] NET38[2] NET38[3] NET37[0]
+NET37[1] NET37[2] NET37[3] NET26[0] NET26[1] NET26[2] NET26[3] NET394 NET393
+NET206 NET389 NET222 NET204 NET32 NET31[0] NET31[1] NET30 NET390 NET231
+NET27[0] NET27[1] NET27[2] NET27[3] NET27[4] NET27[5] NET27[6] NET391[0]
+NET391[1] NET391[2] NET391[3] NET391[4] NET391[5] NET391[6] NET25[0] NET25[1]
+NET25[2] NET25[3] NET392[0] NET392[1] NET392[2] NET392[3] S1100W8_CTRL844_M16
XI10 NET428 NET444 NET479 NET445 NET97 NET96 NET94 NET93 NET92 NET91 NET90[0]
+NET90[1] NET90[2] NET90[3] NET90[4] NET90[5] NET90[6] NET90[7] NET89[0]
+NET89[1] NET89[2] NET89[3] NET88[0] NET88[1] NET88[2] NET88[3] NET87[0]
+NET87[1] NET87[2] NET87[3] NET76[0] NET76[1] NET421 NET420 NET86 NET426 NET85
+NET83 NET82 NET81[0] NET81[1] NET80 NET424 NET235 NET77[0] NET77[1] NET77[2]
+NET77[3] NET77[4] NET77[5] NET77[6] NET423[0] NET423[1] NET423[2] NET423[3]
+NET423[4] NET423[5] NET423[6] NET74[0] NET74[1] NET74[2] NET422[0] NET422[1]
+NET422[2] S1100W8_CTRL844_M8
XI9 NET460 NET236 NET505 NET475 NET143 NET142 NET140 NET139 NET138 NET137
+NET136[0] NET136[1] NET136[2] NET136[3] NET136[4] NET136[5] NET136[6]
+NET136[7] NET135[0] NET135[1] NET135[2] NET135[3] NET134[0] NET134[1]
+NET134[2] NET134[3] NET133[0] NET133[1] NET133[2] NET133[3] NET458 NET457
+NET132 NET453 NET131 NET129 NET128 NET127[0] NET127[1] NET126 NET48 NET84
+NET123[0] NET123[1] NET123[2] NET123[3] NET123[4] NET123[5] NET123[6] NET52[0]
+NET52[1] NET52[2] NET52[3] NET52[4] NET52[5] NET52[6] NET122[0] NET122[1]
+NET456[0] NET456[1] S1100W8_CTRL844_M4
XI16 NET227 NET226 NET225 S1100W8_MDEC_TRK
XI1 NET3[0] NET3[1] NET2[0] NET2[1] NET1[0] NET1[1] S1100W8_CELLX4
D7 GND NET322 NDIO W=1.2U L=1.8U
.ENDS S1100W8_LEAFCELL


**** End of leaf cells

.SUBCKT S1100W8_DECODER TRKBL TIEH WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] 
+ WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] 
+ WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] 
+ WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] 
+ WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] 
+ WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] 
+ WL[1] WL[0] TRKWL WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] 
+ XPD0[2] XPD0[1] XPD0[0] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] 
+ XPD2[1] XPD2[0]
XTIEH TIEH S1100W8_SRAM_TIEH
XDECTRK TRKWL WLPY WLPYB0 S1100W8_MDEC_TRK
MP1 VDD TRKWL TRKBL VDD PCH W=2.1U L=0.07U
XDEC0 WL[1] WL[0] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[0]
+  S1100W8_XDRV
XDEC1 WL[2] WL[3] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[0]
+  S1100W8_XDRV
XDEC2 WL[5] WL[4] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[0]
+  S1100W8_XDRV
XDEC3 WL[6] WL[7] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[0]
+  S1100W8_XDRV
XDEC4 WL[9] WL[8] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[0]
+  S1100W8_XDRV
XDEC5 WL[10] WL[11] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[0]
+  S1100W8_XDRV
XDEC6 WL[13] WL[12] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[0]
+  S1100W8_XDRV
XDEC7 WL[14] WL[15] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[0]
+  S1100W8_XDRV
XDEC8 WL[17] WL[16] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[0]
+  S1100W8_XDRV
XDEC9 WL[18] WL[19] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[0]
+  S1100W8_XDRV
XDEC10 WL[21] WL[20] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[0]
+  S1100W8_XDRV
XDEC11 WL[22] WL[23] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[0]
+  S1100W8_XDRV
XDEC12 WL[25] WL[24] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[0]
+  S1100W8_XDRV
XDEC13 WL[26] WL[27] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[0]
+  S1100W8_XDRV
XDEC14 WL[29] WL[28] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[0]
+  S1100W8_XDRV
XDEC15 WL[30] WL[31] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[0]
+  S1100W8_XDRV
XDEC16 WL[33] WL[32] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[1]
+  S1100W8_XDRV
XDEC17 WL[34] WL[35] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[1]
+  S1100W8_XDRV
XDEC18 WL[37] WL[36] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[1]
+  S1100W8_XDRV
XDEC19 WL[38] WL[39] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[1]
+  S1100W8_XDRV
XDEC20 WL[41] WL[40] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[1]
+  S1100W8_XDRV
XDEC21 WL[42] WL[43] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[1]
+  S1100W8_XDRV
XDEC22 WL[45] WL[44] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[1]
+  S1100W8_XDRV
XDEC23 WL[46] WL[47] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[1]
+  S1100W8_XDRV
XDEC24 WL[49] WL[48] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[1]
+  S1100W8_XDRV
XDEC25 WL[50] WL[51] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[1]
+  S1100W8_XDRV
XDEC26 WL[53] WL[52] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[1]
+  S1100W8_XDRV
XDEC27 WL[54] WL[55] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[1]
+  S1100W8_XDRV
XDEC28 WL[57] WL[56] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[1]
+  S1100W8_XDRV
XDEC29 WL[58] WL[59] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[1]
+  S1100W8_XDRV
XDEC30 WL[61] WL[60] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[1]
+  S1100W8_XDRV
XDEC31 WL[62] WL[63] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[1]
+  S1100W8_XDRV
.ENDS

.SUBCKT S1100W8_TRKCOL TRKBL TIEL TRKBLB TRKWL WL[63] WL[62] WL[61] WL[60] 
+ WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] 
+ WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] 
+ WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] 
+ WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] 
+ WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] 
+ WL[3] WL[2] WL[1] WL[0]
XTRKDUM0 EDG32[1] EDG32[2] TRKBL TIEL WL[1] WL[0] S1100W8_TRKDUMX2
XTRKDUM2 EDG32[2] EDG32[3] TRKBL TIEL WL[3] WL[2] S1100W8_TRKDUMX2
XTRKDUM4 EDG32[3] EDG32[4] TRKBL TIEL WL[5] WL[4] S1100W8_TRKDUMX2
XTRKDUM6 EDG32[4] EDG32[5] TRKBL TIEL WL[7] WL[6] S1100W8_TRKDUMX2
XTRKDUM8 EDG32[5] EDG32[6] TRKBL TIEL WL[9] WL[8] S1100W8_TRKDUMX2
XTRKDUM10 EDG32[6] EDG32[7] TRKBL TIEL WL[11] WL[10] S1100W8_TRKDUMX2
XTRKDUM12 EDG32[7] EDG32[8] TRKBL TIEL WL[13] WL[12] S1100W8_TRKDUMX2
XTRKDUM14 EDG32[8] EDG32[9] TRKBL TIEL WL[15] WL[14] S1100W8_TRKDUMX2
XTRKDUM16 EDG32[9] EDG32[10] TRKBL TIEL WL[17] WL[16] S1100W8_TRKDUMX2
XTRKDUM18 EDG32[10] EDG32[11] TRKBL TIEL WL[19] WL[18] S1100W8_TRKDUMX2
XTRKDUM20 EDG32[11] EDG32[12] TRKBL TIEL WL[21] WL[20] S1100W8_TRKDUMX2
XTRKDUM22 EDG32[12] EDG32[13] TRKBL TIEL WL[23] WL[22] S1100W8_TRKDUMX2
XTRKDUM24 EDG32[13] EDG32[14] TRKBL TIEL WL[25] WL[24] S1100W8_TRKDUMX2
XTRKDUM26 EDG32[14] EDG32[15] TRKBL TIEL WL[27] WL[26] S1100W8_TRKDUMX2
XTRKDUM28 EDG32[15] EDG32[16] TRKBL TIEL WL[29] WL[28] S1100W8_TRKDUMX2
XTRKDUM30 EDG32[16] EDG32[17] TRKBL TIEL WL[31] WL[30] S1100W8_TRKDUMX2
XTRKDUM32 EDG32[17] EDG32[18] TRKBL TIEL WL[33] WL[32] S1100W8_TRKDUMX2
XTRKDUM34 EDG32[18] EDG32[19] TRKBL TIEL WL[35] WL[34] S1100W8_TRKDUMX2
XTRKDUM36 EDG32[19] EDG32[20] TRKBL TIEL WL[37] WL[36] S1100W8_TRKDUMX2
XTRKDUM38 EDG32[20] EDG32[21] TRKBL TIEL WL[39] WL[38] S1100W8_TRKDUMX2
XTRKNOR40 EDG32[21] EDG32[22] TRKBL TRKBLB TRKWL WL[41] WL[40]
+  S1100W8_TRKNORX2
XTRKNOR42 EDG32[22] EDG32[23] TRKBL TRKBLB TRKWL WL[43] WL[42]
+  S1100W8_TRKNORX2
XTRKNOR44 EDG32[23] EDG32[24] TRKBL TRKBLB TRKWL WL[45] WL[44]
+  S1100W8_TRKNORX2
XTRKNOR46 EDG32[24] EDG32[25] TRKBL TRKBLB TRKWL WL[47] WL[46]
+  S1100W8_TRKNORX2
XTRKNOR48 EDG32[25] EDG32[26] TRKBL TRKBLB TRKWL WL[49] WL[48]
+  S1100W8_TRKNORX2
XTRKNOR50 EDG32[26] EDG32[27] TRKBL TRKBLB TRKWL WL[51] WL[50]
+  S1100W8_TRKNORX2
XTRKNOR52 EDG32[27] EDG32[28] TRKBL TRKBLB TRKWL WL[53] WL[52]
+  S1100W8_TRKNORX2
XTRKNOR54 EDG32[28] EDG32[29] TRKBL TRKBLB TRKWL WL[55] WL[54]
+  S1100W8_TRKNORX2
XTRKNOR56 EDG32[29] EDG32[30] TRKBL TRKBLB TRKWL WL[57] WL[56]
+  S1100W8_TRKNORX2
XTRKNOR58 EDG32[30] EDG32[31] TRKBL TRKBLB TRKWL WL[59] WL[58]
+  S1100W8_TRKNORX2
XTRKNOR60 EDG32[31] EDG32[32] TRKBL TRKBLB TRKWL WL[61] WL[60]
+  S1100W8_TRKNORX2
XTRKNOR62 EDG32[32] EDG32[33] TRKBL TRKBLB TRKWL WL[63] WL[62]
+  S1100W8_TRKNORX2
.ENDS

.SUBCKT S1100W8_CORECOLUMN BL0 BL1 BLB0 BLB1 WL[0] WL[1] WL[2] WL[3] WL[4] 
+ WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] 
+ WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] 
+ WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] 
+ WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] 
+ WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] 
+ WL[60] WL[61] WL[62] WL[63]
XBITCELLX2_0 BL0 BL1 BLB0 BLB1 WL[0] WL[1] S1100W8_CELLX4
XBITCELLX2_1 BL0 BL1 BLB0 BLB1 WL[2] WL[3] S1100W8_CELLX4
XBITCELLX2_2 BL0 BL1 BLB0 BLB1 WL[4] WL[5] S1100W8_CELLX4
XBITCELLX2_3 BL0 BL1 BLB0 BLB1 WL[6] WL[7] S1100W8_CELLX4
XBITCELLX2_4 BL0 BL1 BLB0 BLB1 WL[8] WL[9] S1100W8_CELLX4
XBITCELLX2_5 BL0 BL1 BLB0 BLB1 WL[10] WL[11] S1100W8_CELLX4
XBITCELLX2_6 BL0 BL1 BLB0 BLB1 WL[12] WL[13] S1100W8_CELLX4
XBITCELLX2_7 BL0 BL1 BLB0 BLB1 WL[14] WL[15] S1100W8_CELLX4
XBITCELLX2_8 BL0 BL1 BLB0 BLB1 WL[16] WL[17] S1100W8_CELLX4
XBITCELLX2_9 BL0 BL1 BLB0 BLB1 WL[18] WL[19] S1100W8_CELLX4
XBITCELLX2_10 BL0 BL1 BLB0 BLB1 WL[20] WL[21] S1100W8_CELLX4
XBITCELLX2_11 BL0 BL1 BLB0 BLB1 WL[22] WL[23] S1100W8_CELLX4
XBITCELLX2_12 BL0 BL1 BLB0 BLB1 WL[24] WL[25] S1100W8_CELLX4
XBITCELLX2_13 BL0 BL1 BLB0 BLB1 WL[26] WL[27] S1100W8_CELLX4
XBITCELLX2_14 BL0 BL1 BLB0 BLB1 WL[28] WL[29] S1100W8_CELLX4
XBITCELLX2_15 BL0 BL1 BLB0 BLB1 WL[30] WL[31] S1100W8_CELLX4
XBITCELLX2_16 BL0 BL1 BLB0 BLB1 WL[32] WL[33] S1100W8_CELLX4
XBITCELLX2_17 BL0 BL1 BLB0 BLB1 WL[34] WL[35] S1100W8_CELLX4
XBITCELLX2_18 BL0 BL1 BLB0 BLB1 WL[36] WL[37] S1100W8_CELLX4
XBITCELLX2_19 BL0 BL1 BLB0 BLB1 WL[38] WL[39] S1100W8_CELLX4
XBITCELLX2_20 BL0 BL1 BLB0 BLB1 WL[40] WL[41] S1100W8_CELLX4
XBITCELLX2_21 BL0 BL1 BLB0 BLB1 WL[42] WL[43] S1100W8_CELLX4
XBITCELLX2_22 BL0 BL1 BLB0 BLB1 WL[44] WL[45] S1100W8_CELLX4
XBITCELLX2_23 BL0 BL1 BLB0 BLB1 WL[46] WL[47] S1100W8_CELLX4
XBITCELLX2_24 BL0 BL1 BLB0 BLB1 WL[48] WL[49] S1100W8_CELLX4
XBITCELLX2_25 BL0 BL1 BLB0 BLB1 WL[50] WL[51] S1100W8_CELLX4
XBITCELLX2_26 BL0 BL1 BLB0 BLB1 WL[52] WL[53] S1100W8_CELLX4
XBITCELLX2_27 BL0 BL1 BLB0 BLB1 WL[54] WL[55] S1100W8_CELLX4
XBITCELLX2_28 BL0 BL1 BLB0 BLB1 WL[56] WL[57] S1100W8_CELLX4
XBITCELLX2_29 BL0 BL1 BLB0 BLB1 WL[58] WL[59] S1100W8_CELLX4
XBITCELLX2_30 BL0 BL1 BLB0 BLB1 WL[60] WL[61] S1100W8_CELLX4
XBITCELLX2_31 BL0 BL1 BLB0 BLB1 WL[62] WL[63] S1100W8_CELLX4
.ENDS

.SUBCKT TS1N65LPA256X8M4 Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] A[0] A[1] 
+ A[2] A[3] A[4] A[5] A[6] A[7] BWEB[0] BWEB[1] BWEB[2] BWEB[3] BWEB[4] BWEB[5] 
+ BWEB[6] BWEB[7] CEB CLK D[0] D[1] D[2] D[3] D[4] D[5] D[6] D[7] WEB TSEL[0] 
+ TSEL[1]
XLCOLUMN0 BL[0] BL[1] BLB[0] BLB[1] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN1 BL[2] BL[3] BLB[2] BLB[3] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN2 BL[4] BL[5] BLB[4] BLB[5] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN3 BL[6] BL[7] BLB[6] BLB[7] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN4 BL[8] BL[9] BLB[8] BLB[9] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN5 BL[10] BL[11] BLB[10] BLB[11] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN6 BL[12] BL[13] BLB[12] BLB[13] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN7 BL[14] BL[15] BLB[14] BLB[15] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN8 BL[16] BL[17] BLB[16] BLB[17] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN9 BL[18] BL[19] BLB[18] BLB[19] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN10 BL[20] BL[21] BLB[20] BLB[21] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN11 BL[22] BL[23] BLB[22] BLB[23] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN12 BL[24] BL[25] BLB[24] BLB[25] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN13 BL[26] BL[27] BLB[26] BLB[27] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN14 BL[28] BL[29] BLB[28] BLB[29] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XLCOLUMN15 BL[30] BL[31] BLB[30] BLB[31] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] S1100W8_CORECOLUMN
XIO0 Q[0] BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] AWTI BIST_BUF 
+ BWEB[0] TIELB D[0] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0]
+  S1100W8_IO_M4
XIO1 Q[1] BL[4] BL[5] BL[6] BL[7] BLB[4] BLB[5] BLB[6] BLB[7] AWTI BIST_BUF 
+ BWEB[1] TIELB D[1] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0]
+  S1100W8_IO_M4
XIO2 Q[2] BL[8] BL[9] BL[10] BL[11] BLB[8] BLB[9] BLB[10] BLB[11] AWTI 
+ BIST_BUF BWEB[2] TIELB D[2] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0]
+  S1100W8_IO_M4
XIO3 Q[3] BL[12] BL[13] BL[14] BL[15] BLB[12] BLB[13] BLB[14] BLB[15] AWTI 
+ BIST_BUF BWEB[3] TIELB D[3] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0]
+  S1100W8_IO_M4
XIO4 Q[4] BL[16] BL[17] BL[18] BL[19] BLB[16] BLB[17] BLB[18] BLB[19] AWTI 
+ BIST_BUF BWEB[4] TIELB D[4] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0]
+  S1100W8_IO_M4
XIO5 Q[5] BL[20] BL[21] BL[22] BL[23] BLB[20] BLB[21] BLB[22] BLB[23] AWTI 
+ BIST_BUF BWEB[5] TIELB D[5] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0]
+  S1100W8_IO_M4
XIO6 Q[6] BL[24] BL[25] BL[26] BL[27] BLB[24] BLB[25] BLB[26] BLB[27] AWTI 
+ BIST_BUF BWEB[6] TIELB D[6] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0]
+  S1100W8_IO_M4
XIO7 Q[7] BL[28] BL[29] BL[30] BL[31] BLB[28] BLB[29] BLB[30] BLB[31] AWTI 
+ BIST_BUF BWEB[7] TIELB D[7] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0]
+  S1100W8_IO_M4
XDEC TRKBL TIEH WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] 
+ WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] 
+ WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] 
+ WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] 
+ WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] 
+ WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] TRKWL WLPY
+ WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+ XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0]
+  S1100W8_DECODER
XTRKCOL TRKBL TIEL TIEH TRKWL WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] 
+ WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] 
+ WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] 
+ WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] 
+ WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] 
+ WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] 
+ WL[0] S1100W8_TRKCOL
XCTRL AWTI BIST_BUF TIEL TIELB DCLK GW_RB WLPX WLPY WLPYB0 WLPYB1 XPD0[7] 
+ XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[3] XPD1[2] 
+ XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2] Y10[1] Y10[0] 
+ TIELB TIELB CEB TIELB CLK TIELB TRKBL TSEL[1] TSEL[0] WEB TIELB TIELB TIELB 
+ A[7] A[6] A[5] A[4] A[3] A[2] TIELB TIELB TIELB TIELB TIELB TIELB TIELB A[1] 
+ A[0] TIELB TIELB S1100W8_CTRL844_M4
D0_0 GND A[0] NDIO 0.1066P
D0_1 GND A[1] NDIO 0.1066P
D0_2 GND A[2] NDIO 0.1066P
D0_3 GND A[3] NDIO 0.1066P
D0_4 GND A[4] NDIO 0.1066P
D0_5 GND A[5] NDIO 0.1066P
D0_6 GND A[6] NDIO 0.1066P
D0_7 GND A[7] NDIO 0.1066P
D1_0 GND D[0] NDIO 0.1066P
D10_0 GND BWEB[0] NDIO 0.1066P
D1_1 GND D[1] NDIO 0.1066P
D10_1 GND BWEB[1] NDIO 0.1066P
D1_2 GND D[2] NDIO 0.1066P
D10_2 GND BWEB[2] NDIO 0.1066P
D1_3 GND D[3] NDIO 0.1066P
D10_3 GND BWEB[3] NDIO 0.1066P
D1_4 GND D[4] NDIO 0.1066P
D10_4 GND BWEB[4] NDIO 0.1066P
D1_5 GND D[5] NDIO 0.1066P
D10_5 GND BWEB[5] NDIO 0.1066P
D1_6 GND D[6] NDIO 0.1066P
D10_6 GND BWEB[6] NDIO 0.1066P
D1_7 GND D[7] NDIO 0.1066P
D10_7 GND BWEB[7] NDIO 0.1066P
D2_CEB GND CEB NDIO 0.1066P
D3 GND CLK NDIO 0.1066P
D5 GND WEB NDIO 0.1066P
D9_0 GND TSEL[0] NDIO 0.1066P
D9_1 GND TSEL[1] NDIO 0.1066P
.ENDS


# Created by MC2 : Version 2006.09.01.d on 2024/04/08, 13:51:32

###############################################################################
#        Software       : TSMC MEMORY COMPILER 2006.09.01.d
#        Technology     : 65 nm CMOS LOGIC Low Power LowK Cu 1P9M 1.2
#                         Mix-vt logic, High-vt SRAM
#        Memory Type    : TSMC 65nm low power SP SRAM Without Redundancy
#        Library Name   : ts1n65lpa8192x8m16
#        Library Version: 140a
#        Generated Time : 2024/04/08, 13:51:24
###############################################################################
#
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
#
###############################################################################
 
MACRO TS1N65LPA8192X8M16
	CLASS BLOCK ;
	FOREIGN TS1N65LPA8192X8M16 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 192.940 BY 290.485 ;
	SYMMETRY X Y R90 ;

	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 99.335 0.000 99.855 0.520 ;
			LAYER M2 ;
			RECT 99.335 0.000 99.855 0.520 ;
			LAYER M3 ;
			RECT 99.335 0.000 99.855 0.520 ;
		END
	END A[0]

	PIN A[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 76.675 0.000 77.195 0.520 ;
			LAYER M1 ;
			RECT 76.675 0.000 77.195 0.520 ;
			LAYER M2 ;
			RECT 76.675 0.000 77.195 0.520 ;
		END
	END A[10]

	PIN A[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 73.500 0.000 74.020 0.520 ;
			LAYER M2 ;
			RECT 73.500 0.000 74.020 0.520 ;
			LAYER M3 ;
			RECT 73.500 0.000 74.020 0.520 ;
		END
	END A[11]

	PIN A[12]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 72.055 0.000 72.575 0.520 ;
			LAYER M1 ;
			RECT 72.055 0.000 72.575 0.520 ;
			LAYER M3 ;
			RECT 72.055 0.000 72.575 0.520 ;
		END
	END A[12]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 102.790 0.000 103.310 0.520 ;
			LAYER M3 ;
			RECT 102.790 0.000 103.310 0.520 ;
			LAYER M1 ;
			RECT 102.790 0.000 103.310 0.520 ;
		END
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 103.510 0.000 104.030 0.520 ;
			LAYER M2 ;
			RECT 103.510 0.000 104.030 0.520 ;
			LAYER M3 ;
			RECT 103.510 0.000 104.030 0.520 ;
		END
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 105.670 0.000 106.190 0.520 ;
			LAYER M3 ;
			RECT 105.670 0.000 106.190 0.520 ;
			LAYER M2 ;
			RECT 105.670 0.000 106.190 0.520 ;
		END
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 95.155 0.000 95.675 0.520 ;
			LAYER M3 ;
			RECT 95.155 0.000 95.675 0.520 ;
			LAYER M1 ;
			RECT 95.155 0.000 95.675 0.520 ;
		END
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 91.980 0.000 92.500 0.520 ;
			LAYER M2 ;
			RECT 91.980 0.000 92.500 0.520 ;
			LAYER M1 ;
			RECT 91.980 0.000 92.500 0.520 ;
		END
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 90.535 0.000 91.055 0.520 ;
			LAYER M3 ;
			RECT 90.535 0.000 91.055 0.520 ;
			LAYER M1 ;
			RECT 90.535 0.000 91.055 0.520 ;
		END
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 85.915 0.000 86.435 0.520 ;
			LAYER M2 ;
			RECT 85.915 0.000 86.435 0.520 ;
			LAYER M1 ;
			RECT 85.915 0.000 86.435 0.520 ;
		END
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 82.740 0.000 83.260 0.520 ;
			LAYER M2 ;
			RECT 82.740 0.000 83.260 0.520 ;
			LAYER M3 ;
			RECT 82.740 0.000 83.260 0.520 ;
		END
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 81.295 0.000 81.815 0.520 ;
			LAYER M1 ;
			RECT 81.295 0.000 81.815 0.520 ;
			LAYER M2 ;
			RECT 81.295 0.000 81.815 0.520 ;
		END
	END A[9]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 4.335 0.000 4.855 0.520 ;
			LAYER M2 ;
			RECT 4.335 0.000 4.855 0.520 ;
			LAYER M3 ;
			RECT 4.335 0.000 4.855 0.520 ;
		END
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 21.135 0.000 21.655 0.520 ;
			LAYER M1 ;
			RECT 21.135 0.000 21.655 0.520 ;
			LAYER M2 ;
			RECT 21.135 0.000 21.655 0.520 ;
		END
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 37.935 0.000 38.455 0.520 ;
			LAYER M2 ;
			RECT 37.935 0.000 38.455 0.520 ;
			LAYER M3 ;
			RECT 37.935 0.000 38.455 0.520 ;
		END
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 54.735 0.000 55.255 0.520 ;
			LAYER M1 ;
			RECT 54.735 0.000 55.255 0.520 ;
			LAYER M2 ;
			RECT 54.735 0.000 55.255 0.520 ;
		END
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 137.685 0.000 138.205 0.520 ;
			LAYER M1 ;
			RECT 137.685 0.000 138.205 0.520 ;
			LAYER M2 ;
			RECT 137.685 0.000 138.205 0.520 ;
		END
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 154.485 0.000 155.005 0.520 ;
			LAYER M2 ;
			RECT 154.485 0.000 155.005 0.520 ;
			LAYER M3 ;
			RECT 154.485 0.000 155.005 0.520 ;
		END
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 171.285 0.000 171.805 0.520 ;
			LAYER M1 ;
			RECT 171.285 0.000 171.805 0.520 ;
			LAYER M3 ;
			RECT 171.285 0.000 171.805 0.520 ;
		END
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 188.085 0.000 188.605 0.520 ;
			LAYER M3 ;
			RECT 188.085 0.000 188.605 0.520 ;
			LAYER M1 ;
			RECT 188.085 0.000 188.605 0.520 ;
		END
	END BWEB[7]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 106.390 0.000 106.910 0.520 ;
			LAYER M1 ;
			RECT 106.390 0.000 106.910 0.520 ;
			LAYER M3 ;
			RECT 106.390 0.000 106.910 0.520 ;
		END
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 111.595 0.000 112.115 0.520 ;
			LAYER M1 ;
			RECT 111.595 0.000 112.115 0.520 ;
			LAYER M2 ;
			RECT 111.595 0.000 112.115 0.520 ;
		END
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 2.585 0.000 3.105 0.520 ;
			LAYER M3 ;
			RECT 2.585 0.000 3.105 0.520 ;
			LAYER M2 ;
			RECT 2.585 0.000 3.105 0.520 ;
		END
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 19.385 0.000 19.905 0.520 ;
			LAYER M1 ;
			RECT 19.385 0.000 19.905 0.520 ;
			LAYER M2 ;
			RECT 19.385 0.000 19.905 0.520 ;
		END
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 36.185 0.000 36.705 0.520 ;
			LAYER M3 ;
			RECT 36.185 0.000 36.705 0.520 ;
			LAYER M1 ;
			RECT 36.185 0.000 36.705 0.520 ;
		END
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 52.985 0.000 53.505 0.520 ;
			LAYER M3 ;
			RECT 52.985 0.000 53.505 0.520 ;
			LAYER M1 ;
			RECT 52.985 0.000 53.505 0.520 ;
		END
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 139.435 0.000 139.955 0.520 ;
			LAYER M1 ;
			RECT 139.435 0.000 139.955 0.520 ;
			LAYER M2 ;
			RECT 139.435 0.000 139.955 0.520 ;
		END
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 156.235 0.000 156.755 0.520 ;
			LAYER M2 ;
			RECT 156.235 0.000 156.755 0.520 ;
			LAYER M3 ;
			RECT 156.235 0.000 156.755 0.520 ;
		END
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 173.035 0.000 173.555 0.520 ;
			LAYER M3 ;
			RECT 173.035 0.000 173.555 0.520 ;
			LAYER M1 ;
			RECT 173.035 0.000 173.555 0.520 ;
		END
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 189.835 0.000 190.355 0.520 ;
			LAYER M1 ;
			RECT 189.835 0.000 190.355 0.520 ;
			LAYER M2 ;
			RECT 189.835 0.000 190.355 0.520 ;
		END
	END D[7]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 17.790 0.000 18.310 0.520 ;
			LAYER M1 ;
			RECT 17.790 0.000 18.310 0.520 ;
			LAYER M2 ;
			RECT 17.790 0.000 18.310 0.520 ;
		END
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 34.590 0.000 35.110 0.520 ;
			LAYER M3 ;
			RECT 34.590 0.000 35.110 0.520 ;
			LAYER M1 ;
			RECT 34.590 0.000 35.110 0.520 ;
		END
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 51.390 0.000 51.910 0.520 ;
			LAYER M2 ;
			RECT 51.390 0.000 51.910 0.520 ;
			LAYER M1 ;
			RECT 51.390 0.000 51.910 0.520 ;
		END
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 68.190 0.000 68.710 0.520 ;
			LAYER M1 ;
			RECT 68.190 0.000 68.710 0.520 ;
			LAYER M3 ;
			RECT 68.190 0.000 68.710 0.520 ;
		END
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 124.230 0.000 124.750 0.520 ;
			LAYER M3 ;
			RECT 124.230 0.000 124.750 0.520 ;
			LAYER M1 ;
			RECT 124.230 0.000 124.750 0.520 ;
		END
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 141.030 0.000 141.550 0.520 ;
			LAYER M1 ;
			RECT 141.030 0.000 141.550 0.520 ;
			LAYER M2 ;
			RECT 141.030 0.000 141.550 0.520 ;
		END
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 157.830 0.000 158.350 0.520 ;
			LAYER M2 ;
			RECT 157.830 0.000 158.350 0.520 ;
			LAYER M3 ;
			RECT 157.830 0.000 158.350 0.520 ;
		END
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 174.630 0.000 175.150 0.520 ;
			LAYER M2 ;
			RECT 174.630 0.000 175.150 0.520 ;
			LAYER M1 ;
			RECT 174.630 0.000 175.150 0.520 ;
		END
	END Q[7]

	PIN TSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 119.210 0.000 119.730 0.520 ;
			LAYER M2 ;
			RECT 119.210 0.000 119.730 0.520 ;
			LAYER M1 ;
			RECT 119.210 0.000 119.730 0.520 ;
		END
	END TSEL[0]

	PIN TSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 119.930 0.000 120.450 0.520 ;
			LAYER M3 ;
			RECT 119.930 0.000 120.450 0.520 ;
			LAYER M1 ;
			RECT 119.930 0.000 120.450 0.520 ;
		END
	END TSEL[1]

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 110.340 0.000 110.860 0.520 ;
			LAYER M1 ;
			RECT 110.340 0.000 110.860 0.520 ;
			LAYER M2 ;
			RECT 110.340 0.000 110.860 0.520 ;
		END
	END WEB
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M5 ;
			RECT 0.000 10.000 101.665 14.000 ;
			LAYER M5 ;
			RECT 113.445 10.000 192.940 14.000 ;
			LAYER M5 ;
			RECT 0.000 26.000 101.665 30.000 ;
			LAYER M5 ;
			RECT 113.445 26.000 192.940 30.000 ;
			LAYER M5 ;
			RECT 0.000 42.000 101.665 46.000 ;
			LAYER M5 ;
			RECT 113.445 42.000 192.940 46.000 ;
			LAYER M5 ;
			RECT 0.000 58.000 101.665 62.000 ;
			LAYER M5 ;
			RECT 113.445 58.000 192.940 62.000 ;
			LAYER M5 ;
			RECT 0.000 74.000 101.665 78.000 ;
			LAYER M5 ;
			RECT 113.445 74.000 192.940 78.000 ;
			LAYER M5 ;
			RECT 0.000 90.000 101.665 94.000 ;
			LAYER M5 ;
			RECT 113.445 90.000 192.940 94.000 ;
			LAYER M5 ;
			RECT 0.000 106.000 101.665 110.000 ;
			LAYER M5 ;
			RECT 113.445 106.000 192.940 110.000 ;
			LAYER M5 ;
			RECT 0.000 122.000 101.665 126.000 ;
			LAYER M5 ;
			RECT 113.445 122.000 192.940 126.000 ;
			LAYER M5 ;
			RECT 0.000 138.000 101.665 142.000 ;
			LAYER M5 ;
			RECT 113.445 138.000 192.940 142.000 ;
			LAYER M5 ;
			RECT 0.000 154.000 101.665 158.000 ;
			LAYER M5 ;
			RECT 113.445 154.000 192.940 158.000 ;
			LAYER M5 ;
			RECT 0.000 170.000 101.665 174.000 ;
			LAYER M5 ;
			RECT 113.445 170.000 192.940 174.000 ;
			LAYER M5 ;
			RECT 0.000 186.000 101.665 190.000 ;
			LAYER M5 ;
			RECT 113.445 186.000 192.940 190.000 ;
			LAYER M5 ;
			RECT 0.000 202.000 101.665 206.000 ;
			LAYER M5 ;
			RECT 113.445 202.000 192.940 206.000 ;
			LAYER M5 ;
			RECT 0.000 218.000 101.665 222.000 ;
			LAYER M5 ;
			RECT 113.445 218.000 192.940 222.000 ;
			LAYER M5 ;
			RECT 0.000 234.000 101.665 238.000 ;
			LAYER M5 ;
			RECT 113.445 234.000 192.940 238.000 ;
			LAYER M5 ;
			RECT 0.000 250.000 101.665 254.000 ;
			LAYER M5 ;
			RECT 113.445 250.000 192.940 254.000 ;
			LAYER M5 ;
			RECT 0.000 266.000 101.665 270.000 ;
			LAYER M5 ;
			RECT 113.445 266.000 192.940 270.000 ;
			LAYER M5 ;
			RECT 0.000 282.000 101.665 286.000 ;
			LAYER M5 ;
			RECT 113.445 282.000 192.940 286.000 ;
		LAYER M4 ;
		RECT 0.140 0.730 0.470 290.485 ;
		LAYER M4 ;
		RECT 1.580 0.730 1.960 290.485 ;
		LAYER M4 ;
		RECT 3.680 0.730 4.060 290.485 ;
		LAYER M4 ;
		RECT 5.780 0.730 6.160 290.485 ;
		LAYER M4 ;
		RECT 7.880 0.730 8.260 290.485 ;
		LAYER M4 ;
		RECT 9.980 0.730 10.360 290.485 ;
		LAYER M4 ;
		RECT 12.080 0.730 12.460 290.485 ;
		LAYER M4 ;
		RECT 14.180 0.730 14.560 290.485 ;
		LAYER M4 ;
		RECT 16.280 0.730 16.660 290.485 ;
		LAYER M4 ;
		RECT 18.380 0.730 18.760 290.485 ;
		LAYER M4 ;
		RECT 20.480 0.730 20.860 290.485 ;
		LAYER M4 ;
		RECT 22.580 0.730 22.960 290.485 ;
		LAYER M4 ;
		RECT 24.680 0.730 25.060 290.485 ;
		LAYER M4 ;
		RECT 26.780 0.730 27.160 290.485 ;
		LAYER M4 ;
		RECT 28.880 0.730 29.260 290.485 ;
		LAYER M4 ;
		RECT 30.980 0.730 31.360 290.485 ;
		LAYER M4 ;
		RECT 33.080 0.730 33.460 290.485 ;
		LAYER M4 ;
		RECT 35.180 0.730 35.560 290.485 ;
		LAYER M4 ;
		RECT 37.280 0.730 37.660 290.485 ;
		LAYER M4 ;
		RECT 39.380 0.730 39.760 290.485 ;
		LAYER M4 ;
		RECT 41.480 0.730 41.860 290.485 ;
		LAYER M4 ;
		RECT 43.580 0.730 43.960 290.485 ;
		LAYER M4 ;
		RECT 45.680 0.730 46.060 290.485 ;
		LAYER M4 ;
		RECT 47.780 0.730 48.160 290.485 ;
		LAYER M4 ;
		RECT 49.880 0.730 50.260 290.485 ;
		LAYER M4 ;
		RECT 51.980 0.730 52.360 290.485 ;
		LAYER M4 ;
		RECT 54.080 0.730 54.460 290.485 ;
		LAYER M4 ;
		RECT 56.180 0.730 56.560 290.485 ;
		LAYER M4 ;
		RECT 58.280 0.730 58.660 290.485 ;
		LAYER M4 ;
		RECT 60.380 0.730 60.760 290.485 ;
		LAYER M4 ;
		RECT 62.480 0.730 62.860 290.485 ;
		LAYER M4 ;
		RECT 64.580 0.730 64.960 290.485 ;
		LAYER M4 ;
		RECT 66.680 0.730 67.060 290.485 ;
		LAYER M4 ;
		RECT 68.780 0.730 69.160 290.485 ;
		LAYER M4 ;
		RECT 77.440 0.730 79.800 290.485 ;
		LAYER M4 ;
		RECT 94.505 0.730 97.505 290.485 ;
		LAYER M4 ;
		RECT 106.005 0.730 108.005 290.485 ;
		LAYER M4 ;
		RECT 113.445 0.730 115.445 290.485 ;
		LAYER M4 ;
		RECT 121.680 0.730 122.060 290.485 ;
		LAYER M4 ;
		RECT 123.780 0.730 124.160 290.485 ;
		LAYER M4 ;
		RECT 125.880 0.730 126.260 290.485 ;
		LAYER M4 ;
		RECT 127.980 0.730 128.360 290.485 ;
		LAYER M4 ;
		RECT 130.080 0.730 130.460 290.485 ;
		LAYER M4 ;
		RECT 132.180 0.730 132.560 290.485 ;
		LAYER M4 ;
		RECT 134.280 0.730 134.660 290.485 ;
		LAYER M4 ;
		RECT 136.380 0.730 136.760 290.485 ;
		LAYER M4 ;
		RECT 138.480 0.730 138.860 290.485 ;
		LAYER M4 ;
		RECT 140.580 0.730 140.960 290.485 ;
		LAYER M4 ;
		RECT 142.680 0.730 143.060 290.485 ;
		LAYER M4 ;
		RECT 144.780 0.730 145.160 290.485 ;
		LAYER M4 ;
		RECT 146.880 0.730 147.260 290.485 ;
		LAYER M4 ;
		RECT 148.980 0.730 149.360 290.485 ;
		LAYER M4 ;
		RECT 151.080 0.730 151.460 290.485 ;
		LAYER M4 ;
		RECT 153.180 0.730 153.560 290.485 ;
		LAYER M4 ;
		RECT 155.280 0.730 155.660 290.485 ;
		LAYER M4 ;
		RECT 157.380 0.730 157.760 290.485 ;
		LAYER M4 ;
		RECT 159.480 0.730 159.860 290.485 ;
		LAYER M4 ;
		RECT 161.580 0.730 161.960 290.485 ;
		LAYER M4 ;
		RECT 163.680 0.730 164.060 290.485 ;
		LAYER M4 ;
		RECT 165.780 0.730 166.160 290.485 ;
		LAYER M4 ;
		RECT 167.880 0.730 168.260 290.485 ;
		LAYER M4 ;
		RECT 169.980 0.730 170.360 290.485 ;
		LAYER M4 ;
		RECT 172.080 0.730 172.460 290.485 ;
		LAYER M4 ;
		RECT 174.180 0.730 174.560 290.485 ;
		LAYER M4 ;
		RECT 176.280 0.730 176.660 290.485 ;
		LAYER M4 ;
		RECT 178.380 0.730 178.760 290.485 ;
		LAYER M4 ;
		RECT 180.480 0.730 180.860 290.485 ;
		LAYER M4 ;
		RECT 182.580 0.730 182.960 290.485 ;
		LAYER M4 ;
		RECT 184.680 0.730 185.060 290.485 ;
		LAYER M4 ;
		RECT 186.780 0.730 187.160 290.485 ;
		LAYER M4 ;
		RECT 188.880 0.730 189.260 290.485 ;
		LAYER M4 ;
		RECT 190.980 0.730 191.360 290.485 ;
		LAYER M4 ;
		RECT 192.470 0.730 192.800 290.485 ;
		END
	END VDD

	PIN GND
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M5 ;
			RECT 0.000 2.000 101.665 6.000 ;
			LAYER M5 ;
			RECT 113.445 2.000 192.940 6.000 ;
			LAYER M5 ;
			RECT 0.000 18.000 101.665 22.000 ;
			LAYER M5 ;
			RECT 113.445 18.000 192.940 22.000 ;
			LAYER M5 ;
			RECT 0.000 34.000 101.665 38.000 ;
			LAYER M5 ;
			RECT 113.445 34.000 192.940 38.000 ;
			LAYER M5 ;
			RECT 0.000 50.000 101.665 54.000 ;
			LAYER M5 ;
			RECT 113.445 50.000 192.940 54.000 ;
			LAYER M5 ;
			RECT 0.000 66.000 101.665 70.000 ;
			LAYER M5 ;
			RECT 113.445 66.000 192.940 70.000 ;
			LAYER M5 ;
			RECT 0.000 82.000 101.665 86.000 ;
			LAYER M5 ;
			RECT 113.445 82.000 192.940 86.000 ;
			LAYER M5 ;
			RECT 0.000 98.000 101.665 102.000 ;
			LAYER M5 ;
			RECT 113.445 98.000 192.940 102.000 ;
			LAYER M5 ;
			RECT 0.000 114.000 101.665 118.000 ;
			LAYER M5 ;
			RECT 113.445 114.000 192.940 118.000 ;
			LAYER M5 ;
			RECT 0.000 130.000 101.665 134.000 ;
			LAYER M5 ;
			RECT 113.445 130.000 192.940 134.000 ;
			LAYER M5 ;
			RECT 0.000 146.000 101.665 150.000 ;
			LAYER M5 ;
			RECT 113.445 146.000 192.940 150.000 ;
			LAYER M5 ;
			RECT 0.000 162.000 101.665 166.000 ;
			LAYER M5 ;
			RECT 113.445 162.000 192.940 166.000 ;
			LAYER M5 ;
			RECT 0.000 178.000 101.665 182.000 ;
			LAYER M5 ;
			RECT 113.445 178.000 192.940 182.000 ;
			LAYER M5 ;
			RECT 0.000 194.000 101.665 198.000 ;
			LAYER M5 ;
			RECT 113.445 194.000 192.940 198.000 ;
			LAYER M5 ;
			RECT 0.000 210.000 101.665 214.000 ;
			LAYER M5 ;
			RECT 113.445 210.000 192.940 214.000 ;
			LAYER M5 ;
			RECT 0.000 226.000 101.665 230.000 ;
			LAYER M5 ;
			RECT 113.445 226.000 192.940 230.000 ;
			LAYER M5 ;
			RECT 0.000 242.000 101.665 246.000 ;
			LAYER M5 ;
			RECT 113.445 242.000 192.940 246.000 ;
			LAYER M5 ;
			RECT 0.000 258.000 101.665 262.000 ;
			LAYER M5 ;
			RECT 113.445 258.000 192.940 262.000 ;
			LAYER M5 ;
			RECT 0.000 274.000 101.665 278.000 ;
			LAYER M5 ;
			RECT 113.445 274.000 192.940 278.000 ;
		LAYER M4 ;
		RECT 1.035 0.730 1.415 290.485 ;
		LAYER M4 ;
		RECT 2.530 0.730 3.110 290.485 ;
		LAYER M4 ;
		RECT 4.630 0.730 5.210 290.485 ;
		LAYER M4 ;
		RECT 6.730 0.730 7.310 290.485 ;
		LAYER M4 ;
		RECT 8.830 0.730 9.410 290.485 ;
		LAYER M4 ;
		RECT 10.930 0.730 11.510 290.485 ;
		LAYER M4 ;
		RECT 13.030 0.730 13.610 290.485 ;
		LAYER M4 ;
		RECT 15.130 0.730 15.710 290.485 ;
		LAYER M4 ;
		RECT 17.230 0.730 17.810 290.485 ;
		LAYER M4 ;
		RECT 19.330 0.730 19.910 290.485 ;
		LAYER M4 ;
		RECT 21.430 0.730 22.010 290.485 ;
		LAYER M4 ;
		RECT 23.530 0.730 24.110 290.485 ;
		LAYER M4 ;
		RECT 25.630 0.730 26.210 290.485 ;
		LAYER M4 ;
		RECT 27.730 0.730 28.310 290.485 ;
		LAYER M4 ;
		RECT 29.830 0.730 30.410 290.485 ;
		LAYER M4 ;
		RECT 31.930 0.730 32.510 290.485 ;
		LAYER M4 ;
		RECT 34.030 0.730 34.610 290.485 ;
		LAYER M4 ;
		RECT 36.130 0.730 36.710 290.485 ;
		LAYER M4 ;
		RECT 38.230 0.730 38.810 290.485 ;
		LAYER M4 ;
		RECT 40.330 0.730 40.910 290.485 ;
		LAYER M4 ;
		RECT 42.430 0.730 43.010 290.485 ;
		LAYER M4 ;
		RECT 44.530 0.730 45.110 290.485 ;
		LAYER M4 ;
		RECT 46.630 0.730 47.210 290.485 ;
		LAYER M4 ;
		RECT 48.730 0.730 49.310 290.485 ;
		LAYER M4 ;
		RECT 50.830 0.730 51.410 290.485 ;
		LAYER M4 ;
		RECT 52.930 0.730 53.510 290.485 ;
		LAYER M4 ;
		RECT 55.030 0.730 55.610 290.485 ;
		LAYER M4 ;
		RECT 57.130 0.730 57.710 290.485 ;
		LAYER M4 ;
		RECT 59.230 0.730 59.810 290.485 ;
		LAYER M4 ;
		RECT 61.330 0.730 61.910 290.485 ;
		LAYER M4 ;
		RECT 63.430 0.730 64.010 290.485 ;
		LAYER M4 ;
		RECT 65.530 0.730 66.110 290.485 ;
		LAYER M4 ;
		RECT 67.630 0.730 68.210 290.485 ;
		LAYER M4 ;
		RECT 69.325 0.730 69.705 290.485 ;
		LAYER M4 ;
		RECT 70.205 0.730 73.300 290.485 ;
		LAYER M4 ;
		RECT 93.605 0.730 94.005 290.485 ;
		LAYER M4 ;
		RECT 98.965 0.730 101.665 290.485 ;
		LAYER M4 ;
		RECT 117.370 0.730 120.570 290.485 ;
		LAYER M4 ;
		RECT 121.135 0.730 121.515 290.485 ;
		LAYER M4 ;
		RECT 122.630 0.730 123.210 290.485 ;
		LAYER M4 ;
		RECT 124.730 0.730 125.310 290.485 ;
		LAYER M4 ;
		RECT 126.830 0.730 127.410 290.485 ;
		LAYER M4 ;
		RECT 128.930 0.730 129.510 290.485 ;
		LAYER M4 ;
		RECT 131.030 0.730 131.610 290.485 ;
		LAYER M4 ;
		RECT 133.130 0.730 133.710 290.485 ;
		LAYER M4 ;
		RECT 135.230 0.730 135.810 290.485 ;
		LAYER M4 ;
		RECT 137.330 0.730 137.910 290.485 ;
		LAYER M4 ;
		RECT 139.430 0.730 140.010 290.485 ;
		LAYER M4 ;
		RECT 141.530 0.730 142.110 290.485 ;
		LAYER M4 ;
		RECT 143.630 0.730 144.210 290.485 ;
		LAYER M4 ;
		RECT 145.730 0.730 146.310 290.485 ;
		LAYER M4 ;
		RECT 147.830 0.730 148.410 290.485 ;
		LAYER M4 ;
		RECT 149.930 0.730 150.510 290.485 ;
		LAYER M4 ;
		RECT 152.030 0.730 152.610 290.485 ;
		LAYER M4 ;
		RECT 154.130 0.730 154.710 290.485 ;
		LAYER M4 ;
		RECT 156.230 0.730 156.810 290.485 ;
		LAYER M4 ;
		RECT 158.330 0.730 158.910 290.485 ;
		LAYER M4 ;
		RECT 160.430 0.730 161.010 290.485 ;
		LAYER M4 ;
		RECT 162.530 0.730 163.110 290.485 ;
		LAYER M4 ;
		RECT 164.630 0.730 165.210 290.485 ;
		LAYER M4 ;
		RECT 166.730 0.730 167.310 290.485 ;
		LAYER M4 ;
		RECT 168.830 0.730 169.410 290.485 ;
		LAYER M4 ;
		RECT 170.930 0.730 171.510 290.485 ;
		LAYER M4 ;
		RECT 173.030 0.730 173.610 290.485 ;
		LAYER M4 ;
		RECT 175.130 0.730 175.710 290.485 ;
		LAYER M4 ;
		RECT 177.230 0.730 177.810 290.485 ;
		LAYER M4 ;
		RECT 179.330 0.730 179.910 290.485 ;
		LAYER M4 ;
		RECT 181.430 0.730 182.010 290.485 ;
		LAYER M4 ;
		RECT 183.530 0.730 184.110 290.485 ;
		LAYER M4 ;
		RECT 185.630 0.730 186.210 290.485 ;
		LAYER M4 ;
		RECT 187.730 0.730 188.310 290.485 ;
		LAYER M4 ;
		RECT 189.830 0.730 190.410 290.485 ;
		LAYER M4 ;
		RECT 191.525 0.730 191.905 290.485 ;
		END
	END GND

	OBS
		# Pmesh blockages
		LAYER M5 ;
		RECT 2.000 10.000 99.665 12.000 ;
		LAYER M5 ;
		RECT 115.445 10.000 190.940 12.000 ;
		LAYER M5 ;
		RECT 2.000 26.000 99.665 28.000 ;
		LAYER M5 ;
		RECT 115.445 26.000 190.940 28.000 ;
		LAYER M5 ;
		RECT 2.000 42.000 99.665 44.000 ;
		LAYER M5 ;
		RECT 115.445 42.000 190.940 44.000 ;
		LAYER M5 ;
		RECT 2.000 58.000 99.665 60.000 ;
		LAYER M5 ;
		RECT 115.445 58.000 190.940 60.000 ;
		LAYER M5 ;
		RECT 2.000 74.000 99.665 76.000 ;
		LAYER M5 ;
		RECT 115.445 74.000 190.940 76.000 ;
		LAYER M5 ;
		RECT 2.000 90.000 99.665 92.000 ;
		LAYER M5 ;
		RECT 115.445 90.000 190.940 92.000 ;
		LAYER M5 ;
		RECT 2.000 106.000 99.665 108.000 ;
		LAYER M5 ;
		RECT 115.445 106.000 190.940 108.000 ;
		LAYER M5 ;
		RECT 2.000 122.000 99.665 124.000 ;
		LAYER M5 ;
		RECT 115.445 122.000 190.940 124.000 ;
		LAYER M5 ;
		RECT 2.000 138.000 99.665 140.000 ;
		LAYER M5 ;
		RECT 115.445 138.000 190.940 140.000 ;
		LAYER M5 ;
		RECT 2.000 154.000 99.665 156.000 ;
		LAYER M5 ;
		RECT 115.445 154.000 190.940 156.000 ;
		LAYER M5 ;
		RECT 2.000 170.000 99.665 172.000 ;
		LAYER M5 ;
		RECT 115.445 170.000 190.940 172.000 ;
		LAYER M5 ;
		RECT 2.000 186.000 99.665 188.000 ;
		LAYER M5 ;
		RECT 115.445 186.000 190.940 188.000 ;
		LAYER M5 ;
		RECT 2.000 202.000 99.665 204.000 ;
		LAYER M5 ;
		RECT 115.445 202.000 190.940 204.000 ;
		LAYER M5 ;
		RECT 2.000 218.000 99.665 220.000 ;
		LAYER M5 ;
		RECT 115.445 218.000 190.940 220.000 ;
		LAYER M5 ;
		RECT 2.000 234.000 99.665 236.000 ;
		LAYER M5 ;
		RECT 115.445 234.000 190.940 236.000 ;
		LAYER M5 ;
		RECT 2.000 250.000 99.665 252.000 ;
		LAYER M5 ;
		RECT 115.445 250.000 190.940 252.000 ;
		LAYER M5 ;
		RECT 2.000 266.000 99.665 268.000 ;
		LAYER M5 ;
		RECT 115.445 266.000 190.940 268.000 ;
		LAYER M5 ;
		RECT 2.000 282.000 99.665 284.000 ;
		LAYER M5 ;
		RECT 115.445 282.000 190.940 284.000 ;
		LAYER M5 ;
		RECT 2.000 2.000 99.665 4.000 ;
		LAYER M5 ;
		RECT 115.445 2.000 190.940 4.000 ;
		LAYER M5 ;
		RECT 2.000 18.000 99.665 20.000 ;
		LAYER M5 ;
		RECT 115.445 18.000 190.940 20.000 ;
		LAYER M5 ;
		RECT 2.000 34.000 99.665 36.000 ;
		LAYER M5 ;
		RECT 115.445 34.000 190.940 36.000 ;
		LAYER M5 ;
		RECT 2.000 50.000 99.665 52.000 ;
		LAYER M5 ;
		RECT 115.445 50.000 190.940 52.000 ;
		LAYER M5 ;
		RECT 2.000 66.000 99.665 68.000 ;
		LAYER M5 ;
		RECT 115.445 66.000 190.940 68.000 ;
		LAYER M5 ;
		RECT 2.000 82.000 99.665 84.000 ;
		LAYER M5 ;
		RECT 115.445 82.000 190.940 84.000 ;
		LAYER M5 ;
		RECT 2.000 98.000 99.665 100.000 ;
		LAYER M5 ;
		RECT 115.445 98.000 190.940 100.000 ;
		LAYER M5 ;
		RECT 2.000 114.000 99.665 116.000 ;
		LAYER M5 ;
		RECT 115.445 114.000 190.940 116.000 ;
		LAYER M5 ;
		RECT 2.000 130.000 99.665 132.000 ;
		LAYER M5 ;
		RECT 115.445 130.000 190.940 132.000 ;
		LAYER M5 ;
		RECT 2.000 146.000 99.665 148.000 ;
		LAYER M5 ;
		RECT 115.445 146.000 190.940 148.000 ;
		LAYER M5 ;
		RECT 2.000 162.000 99.665 164.000 ;
		LAYER M5 ;
		RECT 115.445 162.000 190.940 164.000 ;
		LAYER M5 ;
		RECT 2.000 178.000 99.665 180.000 ;
		LAYER M5 ;
		RECT 115.445 178.000 190.940 180.000 ;
		LAYER M5 ;
		RECT 2.000 194.000 99.665 196.000 ;
		LAYER M5 ;
		RECT 115.445 194.000 190.940 196.000 ;
		LAYER M5 ;
		RECT 2.000 210.000 99.665 212.000 ;
		LAYER M5 ;
		RECT 115.445 210.000 190.940 212.000 ;
		LAYER M5 ;
		RECT 2.000 226.000 99.665 228.000 ;
		LAYER M5 ;
		RECT 115.445 226.000 190.940 228.000 ;
		LAYER M5 ;
		RECT 2.000 242.000 99.665 244.000 ;
		LAYER M5 ;
		RECT 115.445 242.000 190.940 244.000 ;
		LAYER M5 ;
		RECT 2.000 258.000 99.665 260.000 ;
		LAYER M5 ;
		RECT 115.445 258.000 190.940 260.000 ;
		LAYER M5 ;
		RECT 2.000 274.000 99.665 276.000 ;
		LAYER M5 ;
		RECT 115.445 274.000 190.940 276.000 ;

		# Mc2Finalize block inhibit statement blockage
		# Promoted blockages
		LAYER M1 ;
		RECT 190.515 0.000 192.940 0.520 ;
		LAYER M3 ;
		RECT 190.515 0.000 192.940 0.520 ;
		LAYER M2 ;
		RECT 171.965 0.000 172.875 0.520 ;
		LAYER M2 ;
		RECT 190.515 0.000 192.940 0.520 ;
		LAYER M3 ;
		RECT 173.715 0.000 174.470 0.520 ;
		LAYER M2 ;
		RECT 173.715 0.000 174.470 0.520 ;
		LAYER M2 ;
		RECT 38.615 0.000 51.230 0.520 ;
		LAYER M1 ;
		RECT 36.865 0.000 37.775 0.520 ;
		LAYER M3 ;
		RECT 36.865 0.000 37.775 0.520 ;
		LAYER M2 ;
		RECT 36.865 0.000 37.775 0.520 ;
		LAYER M3 ;
		RECT 38.615 0.000 51.230 0.520 ;
		LAYER M1 ;
		RECT 38.615 0.000 51.230 0.520 ;
		LAYER M1 ;
		RECT 52.070 0.000 52.825 0.520 ;
		LAYER M2 ;
		RECT 52.070 0.000 52.825 0.520 ;
		LAYER M1 ;
		RECT 53.665 0.000 54.575 0.520 ;
		LAYER M3 ;
		RECT 52.070 0.000 52.825 0.520 ;
		LAYER M3 ;
		RECT 188.765 0.000 189.675 0.520 ;
		LAYER M3 ;
		RECT 175.310 0.000 187.925 0.520 ;
		LAYER M1 ;
		RECT 173.715 0.000 174.470 0.520 ;
		LAYER M1 ;
		RECT 171.965 0.000 172.875 0.520 ;
		LAYER M2 ;
		RECT 55.415 0.000 68.030 0.520 ;
		LAYER M1 ;
		RECT 55.415 0.000 68.030 0.520 ;
		LAYER M2 ;
		RECT 53.665 0.000 54.575 0.520 ;
		LAYER M3 ;
		RECT 53.665 0.000 54.575 0.520 ;
		LAYER M3 ;
		RECT 55.415 0.000 68.030 0.520 ;
		LAYER M2 ;
		RECT 188.765 0.000 189.675 0.520 ;
		LAYER M1 ;
		RECT 188.765 0.000 189.675 0.520 ;
		LAYER M2 ;
		RECT 175.310 0.000 187.925 0.520 ;
		LAYER M1 ;
		RECT 175.310 0.000 187.925 0.520 ;
		LAYER M4 ;
		RECT 191.360 0.730 191.525 290.485 ;
		LAYER M4 ;
		RECT 121.515 0.730 121.680 290.485 ;
		LAYER M4 ;
		RECT 120.570 0.730 121.135 290.485 ;
		LAYER M1 ;
		RECT 2.425 0.520 192.940 290.485 ;
		LAYER M2 ;
		RECT 2.425 0.520 192.940 290.485 ;
		LAYER M3 ;
		RECT 2.425 0.520 192.940 290.485 ;
		LAYER M3 ;
		RECT 3.265 0.000 4.175 0.520 ;
		LAYER M3 ;
		RECT 171.965 0.000 172.875 0.520 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 192.940 290.485 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 192.940 290.485 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 192.940 290.485 ;
		LAYER M2 ;
		RECT 158.510 0.000 171.125 0.520 ;
		LAYER M3 ;
		RECT 141.710 0.000 154.325 0.520 ;
		LAYER M2 ;
		RECT 155.165 0.000 156.075 0.520 ;
		LAYER M1 ;
		RECT 141.710 0.000 154.325 0.520 ;
		LAYER M2 ;
		RECT 141.710 0.000 154.325 0.520 ;
		LAYER M2 ;
		RECT 120.610 0.000 124.070 0.520 ;
		LAYER M1 ;
		RECT 120.610 0.000 124.070 0.520 ;
		LAYER M1 ;
		RECT 111.020 0.000 111.435 0.520 ;
		LAYER M2 ;
		RECT 111.020 0.000 111.435 0.520 ;
		LAYER M2 ;
		RECT 112.275 0.000 119.050 0.520 ;
		LAYER M2 ;
		RECT 138.365 0.000 139.275 0.520 ;
		LAYER M1 ;
		RECT 107.070 0.000 110.180 0.520 ;
		LAYER M2 ;
		RECT 107.070 0.000 110.180 0.520 ;
		LAYER M1 ;
		RECT 74.180 0.000 76.515 0.520 ;
		LAYER M1 ;
		RECT 81.975 0.000 82.580 0.520 ;
		LAYER M2 ;
		RECT 83.420 0.000 85.755 0.520 ;
		LAYER M1 ;
		RECT 83.420 0.000 85.755 0.520 ;
		LAYER M1 ;
		RECT 158.510 0.000 171.125 0.520 ;
		LAYER M3 ;
		RECT 158.510 0.000 171.125 0.520 ;
		LAYER M3 ;
		RECT 120.610 0.000 124.070 0.520 ;
		LAYER M1 ;
		RECT 140.115 0.000 140.870 0.520 ;
		LAYER M3 ;
		RECT 140.115 0.000 140.870 0.520 ;
		LAYER M2 ;
		RECT 140.115 0.000 140.870 0.520 ;
		LAYER M1 ;
		RECT 156.915 0.000 157.670 0.520 ;
		LAYER M2 ;
		RECT 156.915 0.000 157.670 0.520 ;
		LAYER M3 ;
		RECT 156.915 0.000 157.670 0.520 ;
		LAYER M1 ;
		RECT 155.165 0.000 156.075 0.520 ;
		LAYER M3 ;
		RECT 155.165 0.000 156.075 0.520 ;
		LAYER M1 ;
		RECT 138.365 0.000 139.275 0.520 ;
		LAYER M3 ;
		RECT 138.365 0.000 139.275 0.520 ;
		LAYER M1 ;
		RECT 104.190 0.000 105.510 0.520 ;
		LAYER M3 ;
		RECT 124.910 0.000 137.525 0.520 ;
		LAYER M2 ;
		RECT 124.910 0.000 137.525 0.520 ;
		LAYER M1 ;
		RECT 124.910 0.000 137.525 0.520 ;
		LAYER M1 ;
		RECT 112.275 0.000 119.050 0.520 ;
		LAYER M1 ;
		RECT 68.870 0.000 71.895 0.520 ;
		LAYER M2 ;
		RECT 68.870 0.000 71.895 0.520 ;
		LAYER M3 ;
		RECT 68.870 0.000 71.895 0.520 ;
		LAYER M3 ;
		RECT 112.275 0.000 119.050 0.520 ;
		LAYER M3 ;
		RECT 111.020 0.000 111.435 0.520 ;
		LAYER M3 ;
		RECT 107.070 0.000 110.180 0.520 ;
		LAYER M3 ;
		RECT 104.190 0.000 105.510 0.520 ;
		LAYER M2 ;
		RECT 104.190 0.000 105.510 0.520 ;
		LAYER M2 ;
		RECT 95.835 0.000 99.175 0.520 ;
		LAYER M3 ;
		RECT 95.835 0.000 99.175 0.520 ;
		LAYER M1 ;
		RECT 100.015 0.000 102.630 0.520 ;
		LAYER M2 ;
		RECT 100.015 0.000 102.630 0.520 ;
		LAYER M3 ;
		RECT 100.015 0.000 102.630 0.520 ;
		LAYER M2 ;
		RECT 74.180 0.000 76.515 0.520 ;
		LAYER M2 ;
		RECT 77.355 0.000 81.135 0.520 ;
		LAYER M3 ;
		RECT 77.355 0.000 81.135 0.520 ;
		LAYER M3 ;
		RECT 83.420 0.000 85.755 0.520 ;
		LAYER M2 ;
		RECT 81.975 0.000 82.580 0.520 ;
		LAYER M3 ;
		RECT 81.975 0.000 82.580 0.520 ;
		LAYER M2 ;
		RECT 72.735 0.000 73.340 0.520 ;
		LAYER M3 ;
		RECT 72.735 0.000 73.340 0.520 ;
		LAYER M1 ;
		RECT 72.735 0.000 73.340 0.520 ;
		LAYER M1 ;
		RECT 86.595 0.000 90.375 0.520 ;
		LAYER M3 ;
		RECT 91.215 0.000 91.820 0.520 ;
		LAYER M3 ;
		RECT 92.660 0.000 94.995 0.520 ;
		LAYER M1 ;
		RECT 92.660 0.000 94.995 0.520 ;
		LAYER M3 ;
		RECT 86.595 0.000 90.375 0.520 ;
		LAYER M2 ;
		RECT 86.595 0.000 90.375 0.520 ;
		LAYER M3 ;
		RECT 74.180 0.000 76.515 0.520 ;
		LAYER M1 ;
		RECT 95.835 0.000 99.175 0.520 ;
		LAYER M2 ;
		RECT 92.660 0.000 94.995 0.520 ;
		LAYER M1 ;
		RECT 18.470 0.000 19.225 0.520 ;
		LAYER M3 ;
		RECT 20.065 0.000 20.975 0.520 ;
		LAYER M2 ;
		RECT 20.065 0.000 20.975 0.520 ;
		LAYER M2 ;
		RECT 21.815 0.000 34.430 0.520 ;
		LAYER M1 ;
		RECT 20.065 0.000 20.975 0.520 ;
		LAYER M1 ;
		RECT 77.355 0.000 81.135 0.520 ;
		LAYER M1 ;
		RECT 35.270 0.000 36.025 0.520 ;
		LAYER M3 ;
		RECT 35.270 0.000 36.025 0.520 ;
		LAYER M2 ;
		RECT 35.270 0.000 36.025 0.520 ;
		LAYER M2 ;
		RECT 91.215 0.000 91.820 0.520 ;
		LAYER M1 ;
		RECT 91.215 0.000 91.820 0.520 ;
		LAYER M1 ;
		RECT 21.815 0.000 34.430 0.520 ;
		LAYER M4 ;
		RECT 94.005 0.730 94.505 290.485 ;
		LAYER M4 ;
		RECT 69.160 0.730 69.325 290.485 ;
		LAYER M3 ;
		RECT 5.015 0.000 17.630 0.520 ;
		LAYER M4 ;
		RECT 69.705 0.730 70.205 290.485 ;
		LAYER M1 ;
		RECT 5.015 0.000 17.630 0.520 ;
		LAYER M2 ;
		RECT 5.015 0.000 17.630 0.520 ;
		LAYER M4 ;
		RECT 1.415 0.730 1.580 290.485 ;
		LAYER M2 ;
		RECT 0.000 0.000 2.425 290.485 ;
		LAYER M1 ;
		RECT 3.265 0.000 4.175 0.520 ;
		LAYER M2 ;
		RECT 3.265 0.000 4.175 0.520 ;
		LAYER M3 ;
		RECT 0.000 0.000 2.425 290.485 ;
		LAYER M1 ;
		RECT 0.000 0.000 2.425 290.485 ;
		LAYER M2 ;
		RECT 18.470 0.000 19.225 0.520 ;
		LAYER M3 ;
		RECT 18.470 0.000 19.225 0.520 ;
		LAYER M3 ;
		RECT 21.815 0.000 34.430 0.520 ;
	END
	# End of OBS

END TS1N65LPA8192X8M16

END LIBRARY

# Created by MC2 : Version 2006.09.01.d on 2024/04/08, 13:50:43

###############################################################################
#        Software       : TSMC MEMORY COMPILER 2006.09.01.d
#        Technology     : 65 nm CMOS LOGIC Low Power LowK Cu 1P9M 1.2
#                         Mix-vt logic, High-vt SRAM
#        Memory Type    : TSMC 65nm low power SP SRAM Without Redundancy
#        Library Name   : ts1n65lpa4096x8m8
#        Library Version: 140a
#        Generated Time : 2024/04/08, 13:50:39
###############################################################################
#
#STATEMENT OF USE
#
#This information contains confidential and proprietary information of TSMC.
#No part of this information may be reproduced, transmitted, transcribed,
#stored in a retrieval system, or translated into any human or computer
#language, in any form or by any means, electronic, mechanical, magnetic,
#optical, chemical, manual, or otherwise, without the prior written permission
#of TSMC. This information was prepared for informational purpose and is for
#use by TSMC's customers only. TSMC reserves the right to make changes in the
#information at any time and without notice.
#
###############################################################################
 
MACRO TS1N65LPA4096X8M8
	CLASS BLOCK ;
	FOREIGN TS1N65LPA4096X8M8 0.0 0.0 ;
	ORIGIN 0.0 0.0 ;
	SIZE 116.725 BY 296.985 ;
	SYMMETRY X Y R90 ;

	PIN A[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 62.355 0.000 62.875 0.520 ;
			LAYER M1 ;
			RECT 62.355 0.000 62.875 0.520 ;
			LAYER M2 ;
			RECT 62.355 0.000 62.875 0.520 ;
		END
	END A[0]

	PIN A[10]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 40.615 0.000 41.135 0.520 ;
			LAYER M3 ;
			RECT 40.615 0.000 41.135 0.520 ;
			LAYER M2 ;
			RECT 40.615 0.000 41.135 0.520 ;
		END
	END A[10]

	PIN A[11]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 36.855 0.000 37.375 0.520 ;
			LAYER M1 ;
			RECT 36.855 0.000 37.375 0.520 ;
			LAYER M2 ;
			RECT 36.855 0.000 37.375 0.520 ;
		END
	END A[11]

	PIN A[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 66.230 0.000 66.750 0.520 ;
			LAYER M3 ;
			RECT 66.230 0.000 66.750 0.520 ;
			LAYER M2 ;
			RECT 66.230 0.000 66.750 0.520 ;
		END
	END A[1]

	PIN A[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 70.565 0.000 71.085 0.520 ;
			LAYER M1 ;
			RECT 70.565 0.000 71.085 0.520 ;
			LAYER M2 ;
			RECT 70.565 0.000 71.085 0.520 ;
		END
	END A[2]

	PIN A[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 57.535 0.000 58.055 0.520 ;
			LAYER M2 ;
			RECT 57.535 0.000 58.055 0.520 ;
			LAYER M3 ;
			RECT 57.535 0.000 58.055 0.520 ;
		END
	END A[3]

	PIN A[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 55.655 0.000 56.175 0.520 ;
			LAYER M1 ;
			RECT 55.655 0.000 56.175 0.520 ;
			LAYER M2 ;
			RECT 55.655 0.000 56.175 0.520 ;
		END
	END A[4]

	PIN A[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 51.895 0.000 52.415 0.520 ;
			LAYER M3 ;
			RECT 51.895 0.000 52.415 0.520 ;
			LAYER M1 ;
			RECT 51.895 0.000 52.415 0.520 ;
		END
	END A[5]

	PIN A[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 50.015 0.000 50.535 0.520 ;
			LAYER M3 ;
			RECT 50.015 0.000 50.535 0.520 ;
			LAYER M2 ;
			RECT 50.015 0.000 50.535 0.520 ;
		END
	END A[6]

	PIN A[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 48.135 0.000 48.655 0.520 ;
			LAYER M1 ;
			RECT 48.135 0.000 48.655 0.520 ;
			LAYER M3 ;
			RECT 48.135 0.000 48.655 0.520 ;
		END
	END A[7]

	PIN A[8]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 44.375 0.000 44.895 0.520 ;
			LAYER M1 ;
			RECT 44.375 0.000 44.895 0.520 ;
			LAYER M2 ;
			RECT 44.375 0.000 44.895 0.520 ;
		END
	END A[8]

	PIN A[9]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 42.495 0.000 43.015 0.520 ;
			LAYER M1 ;
			RECT 42.495 0.000 43.015 0.520 ;
			LAYER M2 ;
			RECT 42.495 0.000 43.015 0.520 ;
		END
	END A[9]

	PIN BWEB[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 3.665 0.000 4.185 0.520 ;
			LAYER M2 ;
			RECT 3.665 0.000 4.185 0.520 ;
			LAYER M1 ;
			RECT 3.665 0.000 4.185 0.520 ;
		END
	END BWEB[0]

	PIN BWEB[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 12.065 0.000 12.585 0.520 ;
			LAYER M1 ;
			RECT 12.065 0.000 12.585 0.520 ;
			LAYER M2 ;
			RECT 12.065 0.000 12.585 0.520 ;
		END
	END BWEB[1]

	PIN BWEB[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 20.465 0.000 20.985 0.520 ;
			LAYER M1 ;
			RECT 20.465 0.000 20.985 0.520 ;
			LAYER M2 ;
			RECT 20.465 0.000 20.985 0.520 ;
		END
	END BWEB[2]

	PIN BWEB[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 28.865 0.000 29.385 0.520 ;
			LAYER M2 ;
			RECT 28.865 0.000 29.385 0.520 ;
			LAYER M3 ;
			RECT 28.865 0.000 29.385 0.520 ;
		END
	END BWEB[3]

	PIN BWEB[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 87.340 0.000 87.860 0.520 ;
			LAYER M3 ;
			RECT 87.340 0.000 87.860 0.520 ;
			LAYER M1 ;
			RECT 87.340 0.000 87.860 0.520 ;
		END
	END BWEB[4]

	PIN BWEB[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 95.740 0.000 96.260 0.520 ;
			LAYER M2 ;
			RECT 95.740 0.000 96.260 0.520 ;
			LAYER M3 ;
			RECT 95.740 0.000 96.260 0.520 ;
		END
	END BWEB[5]

	PIN BWEB[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 104.140 0.000 104.660 0.520 ;
			LAYER M1 ;
			RECT 104.140 0.000 104.660 0.520 ;
			LAYER M3 ;
			RECT 104.140 0.000 104.660 0.520 ;
		END
	END BWEB[6]

	PIN BWEB[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 112.540 0.000 113.060 0.520 ;
			LAYER M3 ;
			RECT 112.540 0.000 113.060 0.520 ;
			LAYER M2 ;
			RECT 112.540 0.000 113.060 0.520 ;
		END
	END BWEB[7]

	PIN CEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 72.725 0.000 73.245 0.520 ;
			LAYER M3 ;
			RECT 72.725 0.000 73.245 0.520 ;
			LAYER M2 ;
			RECT 72.725 0.000 73.245 0.520 ;
		END
	END CEB

	PIN CLK
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 67.670 0.000 68.190 0.520 ;
			LAYER M3 ;
			RECT 67.670 0.000 68.190 0.520 ;
			LAYER M1 ;
			RECT 67.670 0.000 68.190 0.520 ;
		END
	END CLK

	PIN D[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 8.890 0.000 9.410 0.520 ;
			LAYER M1 ;
			RECT 8.890 0.000 9.410 0.520 ;
			LAYER M2 ;
			RECT 8.890 0.000 9.410 0.520 ;
		END
	END D[0]

	PIN D[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 17.290 0.000 17.810 0.520 ;
			LAYER M3 ;
			RECT 17.290 0.000 17.810 0.520 ;
			LAYER M2 ;
			RECT 17.290 0.000 17.810 0.520 ;
		END
	END D[1]

	PIN D[2]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 25.690 0.000 26.210 0.520 ;
			LAYER M2 ;
			RECT 25.690 0.000 26.210 0.520 ;
			LAYER M1 ;
			RECT 25.690 0.000 26.210 0.520 ;
		END
	END D[2]

	PIN D[3]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 34.090 0.000 34.610 0.520 ;
			LAYER M2 ;
			RECT 34.090 0.000 34.610 0.520 ;
			LAYER M3 ;
			RECT 34.090 0.000 34.610 0.520 ;
		END
	END D[3]

	PIN D[4]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 82.115 0.000 82.635 0.520 ;
			LAYER M1 ;
			RECT 82.115 0.000 82.635 0.520 ;
			LAYER M3 ;
			RECT 82.115 0.000 82.635 0.520 ;
		END
	END D[4]

	PIN D[5]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 90.515 0.000 91.035 0.520 ;
			LAYER M3 ;
			RECT 90.515 0.000 91.035 0.520 ;
			LAYER M1 ;
			RECT 90.515 0.000 91.035 0.520 ;
		END
	END D[5]

	PIN D[6]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 98.915 0.000 99.435 0.520 ;
			LAYER M1 ;
			RECT 98.915 0.000 99.435 0.520 ;
			LAYER M2 ;
			RECT 98.915 0.000 99.435 0.520 ;
		END
	END D[6]

	PIN D[7]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 107.315 0.000 107.835 0.520 ;
			LAYER M3 ;
			RECT 107.315 0.000 107.835 0.520 ;
			LAYER M1 ;
			RECT 107.315 0.000 107.835 0.520 ;
		END
	END D[7]

	PIN Q[0]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 6.170 0.000 6.690 0.520 ;
			LAYER M2 ;
			RECT 6.170 0.000 6.690 0.520 ;
			LAYER M1 ;
			RECT 6.170 0.000 6.690 0.520 ;
		END
	END Q[0]

	PIN Q[1]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 14.570 0.000 15.090 0.520 ;
			LAYER M3 ;
			RECT 14.570 0.000 15.090 0.520 ;
			LAYER M1 ;
			RECT 14.570 0.000 15.090 0.520 ;
		END
	END Q[1]

	PIN Q[2]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 22.970 0.000 23.490 0.520 ;
			LAYER M3 ;
			RECT 22.970 0.000 23.490 0.520 ;
			LAYER M2 ;
			RECT 22.970 0.000 23.490 0.520 ;
		END
	END Q[2]

	PIN Q[3]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 31.370 0.000 31.890 0.520 ;
			LAYER M2 ;
			RECT 31.370 0.000 31.890 0.520 ;
			LAYER M3 ;
			RECT 31.370 0.000 31.890 0.520 ;
		END
	END Q[3]

	PIN Q[4]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 84.835 0.000 85.355 0.520 ;
			LAYER M1 ;
			RECT 84.835 0.000 85.355 0.520 ;
			LAYER M3 ;
			RECT 84.835 0.000 85.355 0.520 ;
		END
	END Q[4]

	PIN Q[5]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 93.235 0.000 93.755 0.520 ;
			LAYER M2 ;
			RECT 93.235 0.000 93.755 0.520 ;
			LAYER M1 ;
			RECT 93.235 0.000 93.755 0.520 ;
		END
	END Q[5]

	PIN Q[6]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M2 ;
			RECT 101.635 0.000 102.155 0.520 ;
			LAYER M3 ;
			RECT 101.635 0.000 102.155 0.520 ;
			LAYER M1 ;
			RECT 101.635 0.000 102.155 0.520 ;
		END
	END Q[6]

	PIN Q[7]
		DIRECTION OUTPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 110.035 0.000 110.555 0.520 ;
			LAYER M2 ;
			RECT 110.035 0.000 110.555 0.520 ;
			LAYER M1 ;
			RECT 110.035 0.000 110.555 0.520 ;
		END
	END Q[7]

	PIN TSEL[0]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 78.170 0.000 78.690 0.520 ;
			LAYER M2 ;
			RECT 78.170 0.000 78.690 0.520 ;
			LAYER M1 ;
			RECT 78.170 0.000 78.690 0.520 ;
		END
	END TSEL[0]

	PIN TSEL[1]
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M3 ;
			RECT 80.085 0.000 80.605 0.520 ;
			LAYER M1 ;
			RECT 80.085 0.000 80.605 0.520 ;
			LAYER M2 ;
			RECT 80.085 0.000 80.605 0.520 ;
		END
	END TSEL[1]

	PIN WEB
		DIRECTION INPUT ;
		USE SIGNAL ;
		PORT
			LAYER M1 ;
			RECT 73.445 0.000 73.965 0.520 ;
			LAYER M3 ;
			RECT 73.445 0.000 73.965 0.520 ;
			LAYER M2 ;
			RECT 73.445 0.000 73.965 0.520 ;
		END
	END WEB
	PIN VDD
		DIRECTION INOUT ;
		USE POWER ;
		PORT
			LAYER M5 ;
			RECT 0.000 10.000 59.050 14.000 ;
			LAYER M5 ;
			RECT 70.830 10.000 116.725 14.000 ;
			LAYER M5 ;
			RECT 0.000 26.000 59.050 30.000 ;
			LAYER M5 ;
			RECT 70.830 26.000 116.725 30.000 ;
			LAYER M5 ;
			RECT 0.000 42.000 59.050 46.000 ;
			LAYER M5 ;
			RECT 70.830 42.000 116.725 46.000 ;
			LAYER M5 ;
			RECT 0.000 58.000 59.050 62.000 ;
			LAYER M5 ;
			RECT 70.830 58.000 116.725 62.000 ;
			LAYER M5 ;
			RECT 0.000 74.000 59.050 78.000 ;
			LAYER M5 ;
			RECT 70.830 74.000 116.725 78.000 ;
			LAYER M5 ;
			RECT 0.000 90.000 59.050 94.000 ;
			LAYER M5 ;
			RECT 70.830 90.000 116.725 94.000 ;
			LAYER M5 ;
			RECT 0.000 106.000 59.050 110.000 ;
			LAYER M5 ;
			RECT 70.830 106.000 116.725 110.000 ;
			LAYER M5 ;
			RECT 0.000 122.000 59.050 126.000 ;
			LAYER M5 ;
			RECT 70.830 122.000 116.725 126.000 ;
			LAYER M5 ;
			RECT 0.000 138.000 59.050 142.000 ;
			LAYER M5 ;
			RECT 70.830 138.000 116.725 142.000 ;
			LAYER M5 ;
			RECT 0.000 154.000 59.050 158.000 ;
			LAYER M5 ;
			RECT 70.830 154.000 116.725 158.000 ;
			LAYER M5 ;
			RECT 0.000 170.000 59.050 174.000 ;
			LAYER M5 ;
			RECT 70.830 170.000 116.725 174.000 ;
			LAYER M5 ;
			RECT 0.000 186.000 59.050 190.000 ;
			LAYER M5 ;
			RECT 70.830 186.000 116.725 190.000 ;
			LAYER M5 ;
			RECT 0.000 202.000 59.050 206.000 ;
			LAYER M5 ;
			RECT 70.830 202.000 116.725 206.000 ;
			LAYER M5 ;
			RECT 0.000 218.000 59.050 222.000 ;
			LAYER M5 ;
			RECT 70.830 218.000 116.725 222.000 ;
			LAYER M5 ;
			RECT 0.000 234.000 59.050 238.000 ;
			LAYER M5 ;
			RECT 70.830 234.000 116.725 238.000 ;
			LAYER M5 ;
			RECT 0.000 250.000 59.050 254.000 ;
			LAYER M5 ;
			RECT 70.830 250.000 116.725 254.000 ;
			LAYER M5 ;
			RECT 0.000 266.000 59.050 270.000 ;
			LAYER M5 ;
			RECT 70.830 266.000 116.725 270.000 ;
			LAYER M5 ;
			RECT 0.000 282.000 59.050 286.000 ;
			LAYER M5 ;
			RECT 70.830 282.000 116.725 286.000 ;
		LAYER M4 ;
		RECT 0.140 1.000 0.470 296.985 ;
		LAYER M4 ;
		RECT 1.580 1.000 1.960 296.985 ;
		LAYER M4 ;
		RECT 3.680 1.000 4.060 296.985 ;
		LAYER M4 ;
		RECT 5.780 1.000 6.160 296.985 ;
		LAYER M4 ;
		RECT 7.880 1.000 8.260 296.985 ;
		LAYER M4 ;
		RECT 9.980 1.000 10.360 296.985 ;
		LAYER M4 ;
		RECT 12.080 1.000 12.460 296.985 ;
		LAYER M4 ;
		RECT 14.180 1.000 14.560 296.985 ;
		LAYER M4 ;
		RECT 16.280 1.000 16.660 296.985 ;
		LAYER M4 ;
		RECT 18.380 1.000 18.760 296.985 ;
		LAYER M4 ;
		RECT 20.480 1.000 20.860 296.985 ;
		LAYER M4 ;
		RECT 22.580 1.000 22.960 296.985 ;
		LAYER M4 ;
		RECT 24.680 1.000 25.060 296.985 ;
		LAYER M4 ;
		RECT 26.780 1.000 27.160 296.985 ;
		LAYER M4 ;
		RECT 28.880 1.000 29.260 296.985 ;
		LAYER M4 ;
		RECT 30.980 1.000 31.360 296.985 ;
		LAYER M4 ;
		RECT 33.080 1.000 33.460 296.985 ;
		LAYER M4 ;
		RECT 35.180 1.000 35.560 296.985 ;
		LAYER M4 ;
		RECT 51.890 1.000 54.890 296.985 ;
		LAYER M4 ;
		RECT 63.390 1.000 65.390 296.985 ;
		LAYER M4 ;
		RECT 70.830 1.000 72.830 296.985 ;
		LAYER M4 ;
		RECT 79.065 1.000 79.445 296.985 ;
		LAYER M4 ;
		RECT 81.165 1.000 81.545 296.985 ;
		LAYER M4 ;
		RECT 83.265 1.000 83.645 296.985 ;
		LAYER M4 ;
		RECT 85.365 1.000 85.745 296.985 ;
		LAYER M4 ;
		RECT 87.465 1.000 87.845 296.985 ;
		LAYER M4 ;
		RECT 89.565 1.000 89.945 296.985 ;
		LAYER M4 ;
		RECT 91.665 1.000 92.045 296.985 ;
		LAYER M4 ;
		RECT 93.765 1.000 94.145 296.985 ;
		LAYER M4 ;
		RECT 95.865 1.000 96.245 296.985 ;
		LAYER M4 ;
		RECT 97.965 1.000 98.345 296.985 ;
		LAYER M4 ;
		RECT 100.065 1.000 100.445 296.985 ;
		LAYER M4 ;
		RECT 102.165 1.000 102.545 296.985 ;
		LAYER M4 ;
		RECT 104.265 1.000 104.645 296.985 ;
		LAYER M4 ;
		RECT 106.365 1.000 106.745 296.985 ;
		LAYER M4 ;
		RECT 108.465 1.000 108.845 296.985 ;
		LAYER M4 ;
		RECT 110.565 1.000 110.945 296.985 ;
		LAYER M4 ;
		RECT 112.665 1.000 113.045 296.985 ;
		LAYER M4 ;
		RECT 114.765 1.000 115.145 296.985 ;
		LAYER M4 ;
		RECT 116.255 1.000 116.585 296.985 ;
		END
	END VDD

	PIN GND
		DIRECTION INOUT ;
		USE GROUND ;
		PORT
			LAYER M5 ;
			RECT 0.000 2.000 59.050 6.000 ;
			LAYER M5 ;
			RECT 70.830 2.000 116.725 6.000 ;
			LAYER M5 ;
			RECT 0.000 18.000 59.050 22.000 ;
			LAYER M5 ;
			RECT 70.830 18.000 116.725 22.000 ;
			LAYER M5 ;
			RECT 0.000 34.000 59.050 38.000 ;
			LAYER M5 ;
			RECT 70.830 34.000 116.725 38.000 ;
			LAYER M5 ;
			RECT 0.000 50.000 59.050 54.000 ;
			LAYER M5 ;
			RECT 70.830 50.000 116.725 54.000 ;
			LAYER M5 ;
			RECT 0.000 66.000 59.050 70.000 ;
			LAYER M5 ;
			RECT 70.830 66.000 116.725 70.000 ;
			LAYER M5 ;
			RECT 0.000 82.000 59.050 86.000 ;
			LAYER M5 ;
			RECT 70.830 82.000 116.725 86.000 ;
			LAYER M5 ;
			RECT 0.000 98.000 59.050 102.000 ;
			LAYER M5 ;
			RECT 70.830 98.000 116.725 102.000 ;
			LAYER M5 ;
			RECT 0.000 114.000 59.050 118.000 ;
			LAYER M5 ;
			RECT 70.830 114.000 116.725 118.000 ;
			LAYER M5 ;
			RECT 0.000 130.000 59.050 134.000 ;
			LAYER M5 ;
			RECT 70.830 130.000 116.725 134.000 ;
			LAYER M5 ;
			RECT 0.000 146.000 59.050 150.000 ;
			LAYER M5 ;
			RECT 70.830 146.000 116.725 150.000 ;
			LAYER M5 ;
			RECT 0.000 162.000 59.050 166.000 ;
			LAYER M5 ;
			RECT 70.830 162.000 116.725 166.000 ;
			LAYER M5 ;
			RECT 0.000 178.000 59.050 182.000 ;
			LAYER M5 ;
			RECT 70.830 178.000 116.725 182.000 ;
			LAYER M5 ;
			RECT 0.000 194.000 59.050 198.000 ;
			LAYER M5 ;
			RECT 70.830 194.000 116.725 198.000 ;
			LAYER M5 ;
			RECT 0.000 210.000 59.050 214.000 ;
			LAYER M5 ;
			RECT 70.830 210.000 116.725 214.000 ;
			LAYER M5 ;
			RECT 0.000 226.000 59.050 230.000 ;
			LAYER M5 ;
			RECT 70.830 226.000 116.725 230.000 ;
			LAYER M5 ;
			RECT 0.000 242.000 59.050 246.000 ;
			LAYER M5 ;
			RECT 70.830 242.000 116.725 246.000 ;
			LAYER M5 ;
			RECT 0.000 258.000 59.050 262.000 ;
			LAYER M5 ;
			RECT 70.830 258.000 116.725 262.000 ;
			LAYER M5 ;
			RECT 0.000 274.000 59.050 278.000 ;
			LAYER M5 ;
			RECT 70.830 274.000 116.725 278.000 ;
			LAYER M5 ;
			RECT 0.000 290.000 59.050 294.000 ;
			LAYER M5 ;
			RECT 70.830 290.000 116.725 294.000 ;
		LAYER M4 ;
		RECT 1.035 1.000 1.415 296.985 ;
		LAYER M4 ;
		RECT 2.530 1.000 3.110 296.985 ;
		LAYER M4 ;
		RECT 4.630 1.000 5.210 296.985 ;
		LAYER M4 ;
		RECT 6.730 1.000 7.310 296.985 ;
		LAYER M4 ;
		RECT 8.830 1.000 9.410 296.985 ;
		LAYER M4 ;
		RECT 10.930 1.000 11.510 296.985 ;
		LAYER M4 ;
		RECT 13.030 1.000 13.610 296.985 ;
		LAYER M4 ;
		RECT 15.130 1.000 15.710 296.985 ;
		LAYER M4 ;
		RECT 17.230 1.000 17.810 296.985 ;
		LAYER M4 ;
		RECT 19.330 1.000 19.910 296.985 ;
		LAYER M4 ;
		RECT 21.430 1.000 22.010 296.985 ;
		LAYER M4 ;
		RECT 23.530 1.000 24.110 296.985 ;
		LAYER M4 ;
		RECT 25.630 1.000 26.210 296.985 ;
		LAYER M4 ;
		RECT 27.730 1.000 28.310 296.985 ;
		LAYER M4 ;
		RECT 29.830 1.000 30.410 296.985 ;
		LAYER M4 ;
		RECT 31.930 1.000 32.510 296.985 ;
		LAYER M4 ;
		RECT 34.030 1.000 34.610 296.985 ;
		LAYER M4 ;
		RECT 35.725 1.000 36.105 296.985 ;
		LAYER M4 ;
		RECT 36.605 1.000 38.605 296.985 ;
		LAYER M4 ;
		RECT 50.990 1.000 51.390 296.985 ;
		LAYER M4 ;
		RECT 56.350 1.000 59.050 296.985 ;
		LAYER M4 ;
		RECT 74.755 1.000 77.955 296.985 ;
		LAYER M4 ;
		RECT 78.520 1.000 78.900 296.985 ;
		LAYER M4 ;
		RECT 80.015 1.000 80.595 296.985 ;
		LAYER M4 ;
		RECT 82.115 1.000 82.695 296.985 ;
		LAYER M4 ;
		RECT 84.215 1.000 84.795 296.985 ;
		LAYER M4 ;
		RECT 86.315 1.000 86.895 296.985 ;
		LAYER M4 ;
		RECT 88.415 1.000 88.995 296.985 ;
		LAYER M4 ;
		RECT 90.515 1.000 91.095 296.985 ;
		LAYER M4 ;
		RECT 92.615 1.000 93.195 296.985 ;
		LAYER M4 ;
		RECT 94.715 1.000 95.295 296.985 ;
		LAYER M4 ;
		RECT 96.815 1.000 97.395 296.985 ;
		LAYER M4 ;
		RECT 98.915 1.000 99.495 296.985 ;
		LAYER M4 ;
		RECT 101.015 1.000 101.595 296.985 ;
		LAYER M4 ;
		RECT 103.115 1.000 103.695 296.985 ;
		LAYER M4 ;
		RECT 105.215 1.000 105.795 296.985 ;
		LAYER M4 ;
		RECT 107.315 1.000 107.895 296.985 ;
		LAYER M4 ;
		RECT 109.415 1.000 109.995 296.985 ;
		LAYER M4 ;
		RECT 111.515 1.000 112.095 296.985 ;
		LAYER M4 ;
		RECT 113.615 1.000 114.195 296.985 ;
		LAYER M4 ;
		RECT 115.310 1.000 115.690 296.985 ;
		END
	END GND

	OBS
		# Pmesh blockages
		LAYER M5 ;
		RECT 2.000 10.000 57.050 12.000 ;
		LAYER M5 ;
		RECT 72.830 10.000 114.725 12.000 ;
		LAYER M5 ;
		RECT 2.000 26.000 57.050 28.000 ;
		LAYER M5 ;
		RECT 72.830 26.000 114.725 28.000 ;
		LAYER M5 ;
		RECT 2.000 42.000 57.050 44.000 ;
		LAYER M5 ;
		RECT 72.830 42.000 114.725 44.000 ;
		LAYER M5 ;
		RECT 2.000 58.000 57.050 60.000 ;
		LAYER M5 ;
		RECT 72.830 58.000 114.725 60.000 ;
		LAYER M5 ;
		RECT 2.000 74.000 57.050 76.000 ;
		LAYER M5 ;
		RECT 72.830 74.000 114.725 76.000 ;
		LAYER M5 ;
		RECT 2.000 90.000 57.050 92.000 ;
		LAYER M5 ;
		RECT 72.830 90.000 114.725 92.000 ;
		LAYER M5 ;
		RECT 2.000 106.000 57.050 108.000 ;
		LAYER M5 ;
		RECT 72.830 106.000 114.725 108.000 ;
		LAYER M5 ;
		RECT 2.000 122.000 57.050 124.000 ;
		LAYER M5 ;
		RECT 72.830 122.000 114.725 124.000 ;
		LAYER M5 ;
		RECT 2.000 138.000 57.050 140.000 ;
		LAYER M5 ;
		RECT 72.830 138.000 114.725 140.000 ;
		LAYER M5 ;
		RECT 2.000 154.000 57.050 156.000 ;
		LAYER M5 ;
		RECT 72.830 154.000 114.725 156.000 ;
		LAYER M5 ;
		RECT 2.000 170.000 57.050 172.000 ;
		LAYER M5 ;
		RECT 72.830 170.000 114.725 172.000 ;
		LAYER M5 ;
		RECT 2.000 186.000 57.050 188.000 ;
		LAYER M5 ;
		RECT 72.830 186.000 114.725 188.000 ;
		LAYER M5 ;
		RECT 2.000 202.000 57.050 204.000 ;
		LAYER M5 ;
		RECT 72.830 202.000 114.725 204.000 ;
		LAYER M5 ;
		RECT 2.000 218.000 57.050 220.000 ;
		LAYER M5 ;
		RECT 72.830 218.000 114.725 220.000 ;
		LAYER M5 ;
		RECT 2.000 234.000 57.050 236.000 ;
		LAYER M5 ;
		RECT 72.830 234.000 114.725 236.000 ;
		LAYER M5 ;
		RECT 2.000 250.000 57.050 252.000 ;
		LAYER M5 ;
		RECT 72.830 250.000 114.725 252.000 ;
		LAYER M5 ;
		RECT 2.000 266.000 57.050 268.000 ;
		LAYER M5 ;
		RECT 72.830 266.000 114.725 268.000 ;
		LAYER M5 ;
		RECT 2.000 282.000 57.050 284.000 ;
		LAYER M5 ;
		RECT 72.830 282.000 114.725 284.000 ;
		LAYER M5 ;
		RECT 2.000 2.000 57.050 4.000 ;
		LAYER M5 ;
		RECT 72.830 2.000 114.725 4.000 ;
		LAYER M5 ;
		RECT 2.000 18.000 57.050 20.000 ;
		LAYER M5 ;
		RECT 72.830 18.000 114.725 20.000 ;
		LAYER M5 ;
		RECT 2.000 34.000 57.050 36.000 ;
		LAYER M5 ;
		RECT 72.830 34.000 114.725 36.000 ;
		LAYER M5 ;
		RECT 2.000 50.000 57.050 52.000 ;
		LAYER M5 ;
		RECT 72.830 50.000 114.725 52.000 ;
		LAYER M5 ;
		RECT 2.000 66.000 57.050 68.000 ;
		LAYER M5 ;
		RECT 72.830 66.000 114.725 68.000 ;
		LAYER M5 ;
		RECT 2.000 82.000 57.050 84.000 ;
		LAYER M5 ;
		RECT 72.830 82.000 114.725 84.000 ;
		LAYER M5 ;
		RECT 2.000 98.000 57.050 100.000 ;
		LAYER M5 ;
		RECT 72.830 98.000 114.725 100.000 ;
		LAYER M5 ;
		RECT 2.000 114.000 57.050 116.000 ;
		LAYER M5 ;
		RECT 72.830 114.000 114.725 116.000 ;
		LAYER M5 ;
		RECT 2.000 130.000 57.050 132.000 ;
		LAYER M5 ;
		RECT 72.830 130.000 114.725 132.000 ;
		LAYER M5 ;
		RECT 2.000 146.000 57.050 148.000 ;
		LAYER M5 ;
		RECT 72.830 146.000 114.725 148.000 ;
		LAYER M5 ;
		RECT 2.000 162.000 57.050 164.000 ;
		LAYER M5 ;
		RECT 72.830 162.000 114.725 164.000 ;
		LAYER M5 ;
		RECT 2.000 178.000 57.050 180.000 ;
		LAYER M5 ;
		RECT 72.830 178.000 114.725 180.000 ;
		LAYER M5 ;
		RECT 2.000 194.000 57.050 196.000 ;
		LAYER M5 ;
		RECT 72.830 194.000 114.725 196.000 ;
		LAYER M5 ;
		RECT 2.000 210.000 57.050 212.000 ;
		LAYER M5 ;
		RECT 72.830 210.000 114.725 212.000 ;
		LAYER M5 ;
		RECT 2.000 226.000 57.050 228.000 ;
		LAYER M5 ;
		RECT 72.830 226.000 114.725 228.000 ;
		LAYER M5 ;
		RECT 2.000 242.000 57.050 244.000 ;
		LAYER M5 ;
		RECT 72.830 242.000 114.725 244.000 ;
		LAYER M5 ;
		RECT 2.000 258.000 57.050 260.000 ;
		LAYER M5 ;
		RECT 72.830 258.000 114.725 260.000 ;
		LAYER M5 ;
		RECT 2.000 274.000 57.050 276.000 ;
		LAYER M5 ;
		RECT 72.830 274.000 114.725 276.000 ;
		LAYER M5 ;
		RECT 2.000 290.000 57.050 292.000 ;
		LAYER M5 ;
		RECT 72.830 290.000 114.725 292.000 ;

		# Mc2Finalize block inhibit statement blockage
		# Promoted blockages
		LAYER M4 ;
		RECT 115.145 1.000 115.310 296.985 ;
		LAYER M2 ;
		RECT 110.715 0.000 112.380 0.520 ;
		LAYER M3 ;
		RECT 110.715 0.000 112.380 0.520 ;
		LAYER M1 ;
		RECT 107.995 0.000 109.875 0.520 ;
		LAYER M2 ;
		RECT 107.995 0.000 109.875 0.520 ;
		LAYER M3 ;
		RECT 107.995 0.000 109.875 0.520 ;
		LAYER M1 ;
		RECT 110.715 0.000 112.380 0.520 ;
		LAYER M1 ;
		RECT 102.315 0.000 103.980 0.520 ;
		LAYER M1 ;
		RECT 113.220 0.000 116.725 0.520 ;
		LAYER M1 ;
		RECT 104.820 0.000 107.155 0.520 ;
		LAYER M2 ;
		RECT 104.820 0.000 107.155 0.520 ;
		LAYER M3 ;
		RECT 104.820 0.000 107.155 0.520 ;
		LAYER M3 ;
		RECT 113.220 0.000 116.725 0.520 ;
		LAYER M2 ;
		RECT 102.315 0.000 103.980 0.520 ;
		LAYER M3 ;
		RECT 102.315 0.000 103.980 0.520 ;
		LAYER M2 ;
		RECT 113.220 0.000 116.725 0.520 ;
		LAYER M2 ;
		RECT 85.515 0.000 87.180 0.520 ;
		LAYER M3 ;
		RECT 82.795 0.000 84.675 0.520 ;
		LAYER M2 ;
		RECT 82.795 0.000 84.675 0.520 ;
		LAYER M1 ;
		RECT 82.795 0.000 84.675 0.520 ;
		LAYER M1 ;
		RECT 91.195 0.000 93.075 0.520 ;
		LAYER M3 ;
		RECT 88.020 0.000 90.355 0.520 ;
		LAYER M1 ;
		RECT 88.020 0.000 90.355 0.520 ;
		LAYER M2 ;
		RECT 88.020 0.000 90.355 0.520 ;
		LAYER M1 ;
		RECT 99.595 0.000 101.475 0.520 ;
		LAYER M2 ;
		RECT 99.595 0.000 101.475 0.520 ;
		LAYER M3 ;
		RECT 99.595 0.000 101.475 0.520 ;
		LAYER M1 ;
		RECT 96.420 0.000 98.755 0.520 ;
		LAYER M3 ;
		RECT 96.420 0.000 98.755 0.520 ;
		LAYER M2 ;
		RECT 91.195 0.000 93.075 0.520 ;
		LAYER M3 ;
		RECT 91.195 0.000 93.075 0.520 ;
		LAYER M2 ;
		RECT 96.420 0.000 98.755 0.520 ;
		LAYER M3 ;
		RECT 93.915 0.000 95.580 0.520 ;
		LAYER M1 ;
		RECT 93.915 0.000 95.580 0.520 ;
		LAYER M2 ;
		RECT 93.915 0.000 95.580 0.520 ;
		LAYER M1 ;
		RECT 68.350 0.000 70.405 0.520 ;
		LAYER M2 ;
		RECT 68.350 0.000 70.405 0.520 ;
		LAYER M2 ;
		RECT 80.765 0.000 81.955 0.520 ;
		LAYER M3 ;
		RECT 80.765 0.000 81.955 0.520 ;
		LAYER M4 ;
		RECT 1.415 1.000 1.580 296.985 ;
		LAYER M1 ;
		RECT 0.000 0.000 3.505 296.985 ;
		LAYER M4 ;
		RECT 36.105 1.000 36.605 296.985 ;
		LAYER M4 ;
		RECT 35.560 1.000 35.725 296.985 ;
		LAYER M2 ;
		RECT 0.000 0.000 3.505 296.985 ;
		LAYER M3 ;
		RECT 0.000 0.000 3.505 296.985 ;
		LAYER M3 ;
		RECT 85.515 0.000 87.180 0.520 ;
		LAYER M4 ;
		RECT 78.900 1.000 79.065 296.985 ;
		LAYER M4 ;
		RECT 77.955 1.000 78.520 296.985 ;
		LAYER M3 ;
		RECT 63.035 0.000 66.070 0.520 ;
		LAYER VIA3 ;
		RECT 0.000 0.000 116.725 296.985 ;
		LAYER M3 ;
		RECT 3.505 0.520 116.725 296.985 ;
		LAYER VIA2 ;
		RECT 0.000 0.000 116.725 296.985 ;
		LAYER VIA1 ;
		RECT 0.000 0.000 116.725 296.985 ;
		LAYER M3 ;
		RECT 50.695 0.000 51.735 0.520 ;
		LAYER M4 ;
		RECT 51.390 1.000 51.890 296.985 ;
		LAYER M1 ;
		RECT 3.505 0.520 116.725 296.985 ;
		LAYER M2 ;
		RECT 3.505 0.520 116.725 296.985 ;
		LAYER M2 ;
		RECT 41.295 0.000 42.335 0.520 ;
		LAYER M1 ;
		RECT 43.175 0.000 44.215 0.520 ;
		LAYER M3 ;
		RECT 43.175 0.000 44.215 0.520 ;
		LAYER M2 ;
		RECT 45.055 0.000 47.975 0.520 ;
		LAYER M1 ;
		RECT 37.535 0.000 40.455 0.520 ;
		LAYER M1 ;
		RECT 41.295 0.000 42.335 0.520 ;
		LAYER M1 ;
		RECT 34.770 0.000 36.695 0.520 ;
		LAYER M3 ;
		RECT 34.770 0.000 36.695 0.520 ;
		LAYER M2 ;
		RECT 32.050 0.000 33.930 0.520 ;
		LAYER M3 ;
		RECT 32.050 0.000 33.930 0.520 ;
		LAYER M1 ;
		RECT 26.370 0.000 28.705 0.520 ;
		LAYER M2 ;
		RECT 26.370 0.000 28.705 0.520 ;
		LAYER M1 ;
		RECT 29.545 0.000 31.210 0.520 ;
		LAYER M3 ;
		RECT 21.145 0.000 22.810 0.520 ;
		LAYER M1 ;
		RECT 21.145 0.000 22.810 0.520 ;
		LAYER M2 ;
		RECT 21.145 0.000 22.810 0.520 ;
		LAYER M2 ;
		RECT 23.650 0.000 25.530 0.520 ;
		LAYER M2 ;
		RECT 37.535 0.000 40.455 0.520 ;
		LAYER M3 ;
		RECT 37.535 0.000 40.455 0.520 ;
		LAYER M2 ;
		RECT 34.770 0.000 36.695 0.520 ;
		LAYER M1 ;
		RECT 80.765 0.000 81.955 0.520 ;
		LAYER M3 ;
		RECT 66.910 0.000 67.510 0.520 ;
		LAYER M3 ;
		RECT 68.350 0.000 70.405 0.520 ;
		LAYER M3 ;
		RECT 74.125 0.000 78.010 0.520 ;
		LAYER M3 ;
		RECT 52.575 0.000 55.495 0.520 ;
		LAYER M1 ;
		RECT 56.335 0.000 57.375 0.520 ;
		LAYER M3 ;
		RECT 56.335 0.000 57.375 0.520 ;
		LAYER M2 ;
		RECT 56.335 0.000 57.375 0.520 ;
		LAYER M2 ;
		RECT 52.575 0.000 55.495 0.520 ;
		LAYER M1 ;
		RECT 52.575 0.000 55.495 0.520 ;
		LAYER M1 ;
		RECT 50.695 0.000 51.735 0.520 ;
		LAYER M2 ;
		RECT 50.695 0.000 51.735 0.520 ;
		LAYER M1 ;
		RECT 58.215 0.000 62.195 0.520 ;
		LAYER M2 ;
		RECT 58.215 0.000 62.195 0.520 ;
		LAYER M3 ;
		RECT 58.215 0.000 62.195 0.520 ;
		LAYER M2 ;
		RECT 63.035 0.000 66.070 0.520 ;
		LAYER M2 ;
		RECT 71.245 0.000 72.565 0.520 ;
		LAYER M1 ;
		RECT 71.245 0.000 72.565 0.520 ;
		LAYER M3 ;
		RECT 71.245 0.000 72.565 0.520 ;
		LAYER M1 ;
		RECT 74.125 0.000 78.010 0.520 ;
		LAYER M1 ;
		RECT 6.850 0.000 8.730 0.520 ;
		LAYER M3 ;
		RECT 6.850 0.000 8.730 0.520 ;
		LAYER M2 ;
		RECT 9.570 0.000 11.905 0.520 ;
		LAYER M1 ;
		RECT 32.050 0.000 33.930 0.520 ;
		LAYER M2 ;
		RECT 15.250 0.000 17.130 0.520 ;
		LAYER M3 ;
		RECT 15.250 0.000 17.130 0.520 ;
		LAYER M1 ;
		RECT 9.570 0.000 11.905 0.520 ;
		LAYER M3 ;
		RECT 9.570 0.000 11.905 0.520 ;
		LAYER M1 ;
		RECT 85.515 0.000 87.180 0.520 ;
		LAYER M1 ;
		RECT 4.345 0.000 6.010 0.520 ;
		LAYER M2 ;
		RECT 6.850 0.000 8.730 0.520 ;
		LAYER M2 ;
		RECT 4.345 0.000 6.010 0.520 ;
		LAYER M3 ;
		RECT 4.345 0.000 6.010 0.520 ;
		LAYER M2 ;
		RECT 74.125 0.000 78.010 0.520 ;
		LAYER M1 ;
		RECT 78.850 0.000 79.925 0.520 ;
		LAYER M2 ;
		RECT 78.850 0.000 79.925 0.520 ;
		LAYER M3 ;
		RECT 78.850 0.000 79.925 0.520 ;
		LAYER M1 ;
		RECT 66.910 0.000 67.510 0.520 ;
		LAYER M1 ;
		RECT 63.035 0.000 66.070 0.520 ;
		LAYER M2 ;
		RECT 29.545 0.000 31.210 0.520 ;
		LAYER M3 ;
		RECT 29.545 0.000 31.210 0.520 ;
		LAYER M1 ;
		RECT 45.055 0.000 47.975 0.520 ;
		LAYER M2 ;
		RECT 43.175 0.000 44.215 0.520 ;
		LAYER M2 ;
		RECT 66.910 0.000 67.510 0.520 ;
		LAYER M1 ;
		RECT 17.970 0.000 20.305 0.520 ;
		LAYER M3 ;
		RECT 26.370 0.000 28.705 0.520 ;
		LAYER M3 ;
		RECT 23.650 0.000 25.530 0.520 ;
		LAYER M2 ;
		RECT 17.970 0.000 20.305 0.520 ;
		LAYER M3 ;
		RECT 41.295 0.000 42.335 0.520 ;
		LAYER M3 ;
		RECT 48.815 0.000 49.855 0.520 ;
		LAYER M3 ;
		RECT 45.055 0.000 47.975 0.520 ;
		LAYER M1 ;
		RECT 48.815 0.000 49.855 0.520 ;
		LAYER M2 ;
		RECT 48.815 0.000 49.855 0.520 ;
		LAYER M1 ;
		RECT 15.250 0.000 17.130 0.520 ;
		LAYER M3 ;
		RECT 17.970 0.000 20.305 0.520 ;
		LAYER M1 ;
		RECT 23.650 0.000 25.530 0.520 ;
		LAYER M2 ;
		RECT 12.745 0.000 14.410 0.520 ;
		LAYER M1 ;
		RECT 12.745 0.000 14.410 0.520 ;
		LAYER M3 ;
		RECT 12.745 0.000 14.410 0.520 ;
	END
	# End of OBS

END TS1N65LPA4096X8M8

END LIBRARY

**** Created by MC2: Version 2006.09.01.d on 2024/04/08, 13:50:44 

*****************************************************************************
* CDL NETLIST:
* CELL NAME: LEAFCELL
* NETLISTED ON: DEC 15 15:43:47 2005
*****************************************************************************


*****************************************************************************
* GLOBAL NET DECLARATIONS
*****************************************************************************
*.GLOBAL VDD GND


*****************************************************************************
* PIN CONTROL STATEMENT
*****************************************************************************
*.PIN VDD GND


*****************************************************************************
* BIPOLAR DECLARATIONS
*****************************************************************************


*.LDD
*.BIPOLAR 
*.DIOAREA

*.OPTION SCALE=10E-6

*****************************************************************************
* PARAMETER STATEMENT
*****************************************************************************
.PARAM


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRK_DMY                                                            *
* LAST TIME SAVED: OCT 12 13:39:22 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BLTRK_DMY FLOAT TRBL TRWL WL
MN0 BL0_IN NET37 GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NET37 BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 TRBL TRWL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MN3 FLOAT WL NET37 GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 NET37 BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN NET37 VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S11000X8_BLTRK_DMY


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRK_EDG                                                            *
* LAST TIME SAVED: JUN 30 15:24:03 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BLTRK_EDG BL_CONT TRWL
MN0 BL0_IN NET37 GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NET37 BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 BL_CONT TRWL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 NET37 BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN NET37 VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S11000X8_BLTRK_EDG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKDUM                                                               *
* LAST TIME SAVED: OCT 12 13:39:16 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_TRKDUM BL_CONT FLOAT TRBL TIEL WL
XBLTRK FLOAT TRBL TIEL WL S11000X8_BLTRK_DMY
XI14 BL_CONT TIEL S11000X8_BLTRK_EDG
.ENDS S11000X8_TRKDUM


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKDUMX2                                                             *
* LAST TIME SAVED: OCT  4 16:07:09 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_TRKDUMX2 BL_CONT[1] BL_CONT[0] TRBL TIEL WL[1] WL[0]
XI45 BL_CONT[1] NET12 TRBL TIEL WL[1] S11000X8_TRKDUM
XI46 BL_CONT[0] NET12 TRBL TIEL WL[0] S11000X8_TRKDUM
.ENDS S11000X8_TRKDUMX2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRK                                                                *
* LAST TIME SAVED: OCT  4 16:01:28 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BLTRK FLOAT TRBL TRBLB TRWL WL
MN0 BL0_IN TRBLB GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NET42 BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 TRBL TRWL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MN3 FLOAT WL NET42 GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 TRBLB BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN TRBLB VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S11000X8_BLTRK


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRK_EDG2                                                           *
* LAST TIME SAVED: JUN 30 15:51:02 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BLTRK_EDG2 BL_CONT BL0_IN NPD2 PPU1 PPU2 TRWL
MN2 BL_CONT TRWL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MN0 BL0_IN TRWL GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NPD2 TRWL GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MP0 PPU2 TRWL VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 PPU1 TRWL VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S11000X8_BLTRK_EDG2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKNOR                                                               *
* LAST TIME SAVED: OCT  4 16:04:22 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_TRKNOR BL_CONT FLOAT TRBL TIEH TRWL WL
XCELTRK FLOAT TRBL TIEH TRWL WL S11000X8_BLTRK
XI18 BL_CONT NET22 NET23 NET20 NET21 TRWL S11000X8_BLTRK_EDG2
.ENDS S11000X8_TRKNOR


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKNORX2                                                             *
* LAST TIME SAVED: JUL  7 17:14:05 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_TRKNORX2 BL_CONT[1] BL_CONT[0] TRBL TIEH TRWL WL[1] WL[0]
XI52 BL_CONT[1] NET17 TRBL TIEH TRWL WL[1] S11000X8_TRKNOR
XI51 BL_CONT[0] NET17 TRBL TIEH TRWL WL[0] S11000X8_TRKNOR
.ENDS S11000X8_TRKNORX2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRKMIN                                                             *
* LAST TIME SAVED: MAY 17 15:57:20 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BLTRKMIN TRBL TRBLB TRWL WL
MN0 BL0_IN TRWL GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 NET41 BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 TRBL TRBL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MN3 TRBLB WL NET41 GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 NET41 BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN TRWL VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S11000X8_BLTRKMIN


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BLTRKMIN_EDG                                                         *
* LAST TIME SAVED: JUL  1 10:37:26 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BLTRKMIN_EDG BL_CONT TRBL TRWL
MN0 BL0_IN TRWL GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN1 TRWL BL0_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U 
MN2 BL_CONT TRBL BL0_IN GND NCHPG_HVTSR W=0.09U  L=0.075U
MP0 TRWL BL0_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
MP1 BL0_IN TRWL VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U 
.ENDS S11000X8_BLTRKMIN_EDG


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKMIN                                                               *
* LAST TIME SAVED: OCT 12 14:09:32 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_TRKMIN BL_CONT TRBL TIEH TRWL WL
XTRK_VCCMIN TRBL TIEH TRWL WL S11000X8_BLTRKMIN
XI23 BL_CONT TRBL TRWL S11000X8_BLTRKMIN_EDG
.ENDS S11000X8_TRKMIN


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRKMINX2                                                             *
* LAST TIME SAVED: OCT 12 14:09:24 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_TRKMINX2 BL_CONT[1] BL_CONT[0] TRBL TIEH TRWL WL[1] WL[0]
XI47 BL_CONT[0] TRBL TIEH TRWL WL[0] S11000X8_TRKMIN
XI46 BL_CONT[1] TRBL TIEH TRWL WL[1] S11000X8_TRKMIN
.ENDS S11000X8_TRKMINX2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SINV_HVTP                                                            *
* LAST TIME SAVED: AUG  3 14:45:00 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_SINV_HVTP Y A LN=0.06U WN=0.15U LP=0.06U WP=0.3U
M1 VDD A Y VDD PCH_HVT W=WP L=LP
M0 Y A GND GND NCH W=WN L=LN
.ENDS S11000X8_SINV_HVTP


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SRAM_TIEH                                                            *
* LAST TIME SAVED: OCT 19 14:27:29 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_SRAM_TIEH Z
XI50 Z NET18 S11000X8_SINV_HVTP LN=0.07U WN=2U LP=0.07U WP=8U
MN0 NET18 NET32 GND GND NCH W=0.15U L=0.07U
MP0 VDD NET32 NET32 VDD PCH W=0.3U L=0.07U
MP1 NET32 NET18 VDD VDD PCH W=0.3U L=0.07U
.ENDS S11000X8_SRAM_TIEH


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SINV                                                                 *
* LAST TIME SAVED: APR 15 08:08:15 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_SINV Y A LP=0.06U WP=0.3U LN=0.06U WN=0.15U
M0 Y A GND GND NCH W=WN L=LN
M1 VDD A Y VDD PCH W=WP L=LP
.ENDS S11000X8_SINV


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SNAND3                                                               *
* LAST TIME SAVED: APR 18 16:13:20 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_SNAND3 Y A B C LP3=0.06U WP3=0.3U LP2=0.06U WP2=0.3U LP1=0.06U WP1=0.3U
+LN1=0.06U WN1=0.45U LN2=0.06U WN2=0.45U LN3=0.06U WN3=0.45U
M0 NET14 C GND GND NCH W=WN3 L=LN3
M1 NET17 B NET14 GND NCH W=WN2 L=LN2
M2 Y A NET17 GND NCH W=WN1 L=LN1
M3 VDD A Y VDD PCH W=WP1 L=LP1
M4 VDD B Y VDD PCH W=WP2 L=LP2
M5 VDD C Y VDD PCH W=WP3 L=LP3
.ENDS S11000X8_SNAND3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XDRV                                                                 *
* LAST TIME SAVED: DEC 14 16:50:11 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_XDRV WLOUT[1] WLOUT[0] WLPY WLPYB0 WLPYB1 XPD0 XPD0B XPD1 XPD2
XI288 MWL1 MWL0 S11000X8_SINV LP=0.06U WP=0.8U  LN=0.06U WN=0.8U 
XI295 MWL1A MWL0A S11000X8_SINV LP=0.06U WP=0.8U  LN=0.06U WN=0.8U 
XI296 WLOUT[1] MWL2A S11000X8_SINV_HVTP LN=0.06U WN=5U    LP=0.06U WP=10U    M=2
XI275 WLOUT[0] MWL2 S11000X8_SINV_HVTP LN=0.06U WN=5U    LP=0.06U WP=10U    M=2
MN0 MWL2 MWL1 WLPY GND NCH W=2.0U   L=0.06U
MN1 MWL2A MWL1A WLPY GND NCH W=2.0U   L=0.06U
MP0 VDD MWL1 MWL2 VDD PCH W=2.0U   L=0.06U
MP2 VDD MWL1A MWL2A VDD PCH W=2.0U   L=0.06U
MP3 MWL2A WLPYB0 VDD VDD PCH W=2.0U      L=0.06U
MP1 MWL2 WLPYB1 VDD VDD PCH W=2.0U      L=0.06U
XI290 MWL0A XPD2 XPD1 XPD0B S11000X8_SNAND3 LP3=0.06U WP3=0.15U  LP2=0.06U WP2=0.15U
+LP1=0.06U WP1=0.15U  LN1=0.06U WN1=0.15U  LN2=0.06U WN2=0.15U LN3=0.06U
+WN3=0.15U 
XI282 MWL0 XPD2 XPD1 XPD0 S11000X8_SNAND3 LP3=0.06U WP3=0.15U  LP2=0.06U WP2=0.15U
+LP1=0.06U WP1=0.15U  LN1=0.06U WN1=0.15U  LN2=0.06U WN2=0.15U LN3=0.06U
+WN3=0.15U 
**C2 MWL2 GND 10.372F
**C4 MWL1 GND 3.209F
**C3 MWL0 GND 2.040F
**C5 MWL2A GND 9.991F
**C6 MWL1A GND 3.359F
**C7 MWL0A GND 2.282F
.ENDS S11000X8_XDRV


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XDRVX2                                                               *
* LAST TIME SAVED: JUN 13 11:08:29 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_XDRVX2 WL[3] WL[2] WL[1] WL[0] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2]
+XPD0[1] XPD0[0] XPD1 XPD2
XWLDRV_0 WL[1] WL[0] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1 XPD2 S11000X8_XDRV
XWLDRV_1 WL[2] WL[3] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1 XPD2 S11000X8_XDRV
.ENDS S11000X8_XDRVX2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IOYPASS_M16                                                          *
* LAST TIME SAVED: OCT 12 14:13:51 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IOYPASS_M16 BL BLB DL DLB BLEQB YSEL
*MN0 BL YSEL DL GND NCH W=0.8U L=0.06U
MN0 BL YSEL DL GND NCH W=0.89U L=0.06U
*MN1 BLB YSEL DLB GND NCH W=0.8U L=0.06U
MN1 BLB YSEL DLB GND NCH W=0.89U L=0.06U
MP2 BLB BLEQB BL VDD PCH W=2U L=0.06U
MP0 BL NET47 DL VDD PCH W=0.8U L=0.06U
MP3 VDD BLEQB BLB VDD PCH W=2U L=0.06U
MP1 BLB NET47 DLB VDD PCH W=0.8U L=0.06U
MP4 BL BLEQB VDD VDD PCH W=2U L=0.06U
XI9 NET47 YSEL S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.24U
.ENDS S11000X8_IOYPASS_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DIN                                                                  *
* LAST TIME SAVED: DEC 14 16:50:06 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_DIN AWTD BWEB_M D_M BIST BWEB BWEBM D DM
XI13 BIST_BB BIST_B S11000X8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI12 BIST_B BIST S11000X8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI293 BWEB_M NET16 S11000X8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
XI344 BWC BWT S11000X8_SINV LP=0.15U WP=0.28U LN=0.15U WN=0.15U
XI241 NET14 BWC S11000X8_SINV LP=0.15U WP=0.28U LN=0.15U WN=0.15U
XI242 NET16 NET14 S11000X8_SINV LP=0.1U WP=0.28U LN=0.1U WN=0.15U
XI343 BWT NET107 S11000X8_SINV LP=0.15U WP=0.28U LN=0.15U WN=0.15U
XI85 DT NET110 S11000X8_SINV LP=0.1U WP=0.3U LN=0.1U WN=0.15U
XI83 DC DT S11000X8_SINV LP=0.1U WP=0.3U LN=0.1U WN=0.15U
XI59 D_M NET26 S11000X8_SINV LP=0.07U WP=1.2U LN=0.07U WN=0.6U
XI84 NET26 DC S11000X8_SINV LP=0.2U WP=0.6U LN=0.2U WN=0.3U
**C11 BIST_BB GND 1.596F
**C13 BIST_B GND 1.310F
**C37 NET14 GND 0.680F
**C53 NET16 GND 0.860F
**C23 BWC GND 1.411F
**C14 BWT GND 1.879F
**C12 NET107 GND 1.155F
**C9 DT GND 2.044F
**C2 NET26 GND 1.135F
**C1 DC GND 1.509F
**C10 NET110 GND 1.392F
MP9 NET51 DC AWTD VDD PCH W=0.42U L=0.07U
MP8 VDD BWT NET51 VDD PCH W=0.42U L=0.07U
MP5 VDD BWC NET59 VDD PCH W=0.42U L=0.07U
MP4 NET59 DT AWTD VDD PCH W=0.42U L=0.07U
MP3 NET62 BIST_B NET107 VDD PCH W=0.3U L=0.06U
MP7 VDD BWEBM NET62 VDD PCH W=0.3U L=0.06U
MP1 VDD BWEB NET71 VDD PCH W=0.3U L=0.06U
MP0 NET71 BIST_BB NET107 VDD PCH W=0.3U L=0.06U
MP15 NET74 BIST_BB NET110 VDD PCH W=0.3U L=0.06U
MP14 VDD D NET74 VDD PCH W=0.3U L=0.06U
MP2 VDD DM NET83 VDD PCH W=0.3U L=0.06U
MP6 NET83 BIST_B NET110 VDD PCH W=0.3U L=0.06U
MN7 NET86 BWT GND GND NCH W=0.21U L=0.07U
MN5 AWTD BWC NET86 GND NCH W=0.21U L=0.07U
MN4 AWTD DT NET86 GND NCH W=0.21U L=0.07U
MN3 NET86 DC GND GND NCH W=0.21U L=0.07U
MN6 NET98 BWEBM GND GND NCH W=0.15U L=0.06U
MN2 NET101 BWEB GND GND NCH W=0.15U L=0.06U
MN1 NET107 BIST_BB NET98 GND NCH W=0.15U L=0.06U
MN0 NET107 BIST_B NET101 GND NCH W=0.15U L=0.06U
MN15 NET110 BIST_B NET116 GND NCH W=0.15U L=0.06U
MN14 NET110 BIST_BB NET119 GND NCH W=0.15U L=0.06U
MN13 NET116 D GND GND NCH W=0.15U L=0.06U
MN9 NET119 DM GND GND NCH W=0.15U L=0.06U
.ENDS S11000X8_DIN


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SNOR                                                                 *
* LAST TIME SAVED: APR 15 09:10:54 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_SNOR Y A B LP1=0.06U WP1=0.6U LP2=0.06U WP2=0.6U LN2=0.06U WN2=0.15U LN1=0.06U
+WN1=0.15U
M3 Y A GND GND NCH W=WN1 L=LN1
M2 Y B GND GND NCH W=WN2 L=LN2
M1 NET3 B Y VDD PCH W=WP2 L=LP2
M0 VDD A NET3 VDD PCH W=WP1 L=LP1
.ENDS S11000X8_SNOR


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SA                                                                   *
* LAST TIME SAVED: DEC 14 16:50:07 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_SA Q AWTD AWTI DL DLB PGB PREB SAE
MN11 Z4 AWTD GND GND NCH W=0.9U L=0.07U M=1
MN10 Z4 AWTT Q_B GND NCH W=0.9U L=0.07U M=1
MN8 Z6 AWTC Q_B GND NCH W=0.9U L=0.07U M=1
MN5 Z6 SOB GND GND NCH W=0.9U L=0.07U M=1
MN2 NS SAE GND GND NCH W=2.0U L=0.08U
MN1 DLB_IN DL_IN NS GND NCH W=2.0U L=0.18U
MN0 NS DLB_IN DL_IN GND NCH W=2.0U L=0.18U
MP14 Q_B AWTT Z5 VDD PCH W=1.8U L=0.07U M=1
MP5 Z3 AWTD VDD VDD PCH W=1.8U L=0.07U M=1
MP9 Q_B AWTC Z3 VDD PCH W=1.8U L=0.07U M=1
MP13 Z5 SOB VDD VDD PCH W=1.8U L=0.07U M=1
MP10 VDD PREB DL_IN VDD PCH W=1.0U L=0.1U
MP11 VDD PREB DLB_IN VDD PCH W=1.0U L=0.1U
MP8 DLB_IN PREB DL_IN VDD PCH W=1.2U L=0.12U
MP3 VDD DL_IN DLB_IN VDD PCH W=1.0U L=0.12U
MP2 DL_IN DLB_IN VDD VDD PCH W=1.0U L=0.12U
MP7 DLB PGB DLB_IN VDD PCH W=1.2U L=0.1U
MP6 DL_IN PGB DL VDD PCH W=1.2U L=0.1U
XI152 SO SOB NET096 S11000X8_SNOR LP1=0.07U WP1=2.4U LP2=0.07U WP2=2.4U LN2=0.07U WN2=0.8U
+LN1=0.07U WN1=0.8U
XI116 SOB SO NET098 S11000X8_SNOR LP1=0.07U WP1=2.4U LP2=0.07U WP2=2.4U LN2=0.07U WN2=0.8U
+LN1=0.07U WN1=0.8U
XI153 NET096 DL_IN S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.38U
XI148 NET098 DLB_IN S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.38U
XI61 AWTC AWTI S11000X8_SINV LP=0.06U WP=0.48U LN=0.06U WN=0.24U
XI62 AWTT AWTC S11000X8_SINV LP=0.06U WP=0.48U LN=0.06U WN=0.24U
XI160 Q Q_B S11000X8_SINV LP=0.07U WP=3.6U LN=0.07U WN=1.8U
**C0 DL_IN GND 4.360F
**C1 DLB_IN GND 4.037F
**C4 SO GND 1.951F
**C15 AWTC GND 1.969F
**C7 NET096 GND 2.576F
**C16 AWTT GND 2.078F
**C9 NET098 GND 2.471F
**C14 SOB GND 3.090F
**C17 Q_B GND 2.798F
.ENDS S11000X8_SA


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: TRANSGATE                                                            *
* LAST TIME SAVED: APR 15 08:43:26 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_TRANSGATE Y A C CB LP=0.06U WP=0.3U LN=0.06U WN=0.15U
*.NOPIN VDD GND
M1 A C Y GND NCH W=WN L=LN
M0 Y CB A VDD PCH W=WP L=LP
.ENDS S11000X8_TRANSGATE


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_DCLK                                                              *
* LAST TIME SAVED: DEC 14 16:50:06 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_LH_DCLK Q CP D
**C2 P2 GND 1.709F
**C0 INCP GND 1.251F
XI26 D P2 CP INCP S11000X8_TRANSGATE LP=0.07U WP=0.5U LN=0.07U WN=0.5U
XI33 Q P2 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI29 INCP CP S11000X8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.3U
MN12 GND Q NET39 GND NCH W=0.15U L=0.07U
MN11 NET39 INCP P2 GND NCH W=0.15U L=0.07U
MP4 NET69 Q VDD VDD PCH W=0.28U L=0.07U
MP5 P2 CP NET69 VDD PCH W=0.28U L=0.07U
.ENDS S11000X8_LH_DCLK


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_WRIN_M16                                                          *
* LAST TIME SAVED: SEP 28 10:50:28 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IO_WRIN_M16 DL DLB D DCLK DLEQB WPG
XLH_DCLK_M8 D1B DCLK D S11000X8_LH_DCLK
MP7 DL DLEQB VDD VDD PCH W=1U L=0.07U
MP8 VDD DLEQB DLB VDD PCH W=1U L=0.07U
MN2 VDD D1 D2B VDD PCH W=2.5U L=0.07U
MN0 VDD D1B D2 VDD PCH W=2.5U L=0.07U
MN5 DLB WPG D2B GND NCH W=2.5U L=0.07U
MN4 D2 WPG DL GND NCH W=2.5U L=0.07U
MN3 D2B D1 GND GND NCH W=5U L=0.07U
MN1 D2 D1B GND GND NCH W=5U L=0.07U
XI69 D1 D1B S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
**C11 D1B GND 4.2F
**C6 D1 GND 2.6F
**C7 D2B GND 4.5F
**C8 D2 GND 4.5F
.ENDS S11000X8_IO_WRIN_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_BWEB                                                              *
* LAST TIME SAVED: DEC 14 16:50:07 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_LH_BWEB Q CP D
MP5 P2 CP NET42 VDD PCH W=0.2U L=0.07U
MP4 NET42 Q VDD VDD PCH W=0.2U L=0.07U
XI26 D P2 CP INCP S11000X8_TRANSGATE LP=0.07U WP=0.5U LN=0.07U WN=0.5U
XI29 INCP CP S11000X8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.2U
XI24 Q P2 S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.4U
MN12 GND Q NET51 GND NCH W=0.2U L=0.07U
MN11 NET51 INCP P2 GND NCH W=0.2U L=0.07U
**C1 P2 GND 1.855F
**C0 INCP GND 1.980F
.ENDS S11000X8_LH_BWEB


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SNAND                                                                *
* LAST TIME SAVED: APR 15 08:59:39 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_SNAND Y A B LP2=0.06U WP2=0.3U LP1=0.06U WP1=0.3U LN1=0.06U WN1=0.3U LN2=0.06U
+WN2=0.3U
M0 NET9 B GND GND NCH W=WN2 L=LN2
M1 Y A NET9 GND NCH W=WN1 L=LN1
M2 VDD A Y VDD PCH W=WP1 L=LP1
M3 VDD B Y VDD PCH W=WP2 L=LP2
.ENDS S11000X8_SNAND


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_RWCTRL_M16                                                        *
* LAST TIME SAVED: OCT  7 14:27:13 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IO_RWCTRL_M16 BLEQB DLEQB DLH PGB PREB SAE WPG BWEB DCLK GW_RB WLP
X_LH_BWEB BWEB_SU DLH BWEB S11000X8_LH_BWEB
XI289 PREB NET0100 NET161 S11000X8_SNOR LP1=0.07U WP1=1.2U LP2=0.07U WP2=1.2U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI288 NET161 WLPCD2 NET163 S11000X8_SNOR LP1=0.07U WP1=0.35U LP2=0.07U WP2=0.35U LN2=0.07U
+WN2=0.3U LN1=0.07U WN1=0.3U
XI249 WPG GW_R NET089 S11000X8_SNOR LP1=0.07U WP1=1.0U LP2=0.07U WP2=1.0U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI133 NET073 WLPCD0 NET_110 GW_R S11000X8_SNAND3 LP3=0.07U WP3=1.75U LP2=0.07U WP2=1.75U
+LP1=0.07U WP1=1.75U LN1=0.07U WN1=1.2U LN2=0.07U WN2=1.2U LN3=0.07U WN3=1.2U
XI250 PGB NET166 GW_R S11000X8_SNAND LP2=0.07U WP2=0.84U LP1=0.07U WP1=0.84U LN1=0.07U
+WN1=0.7U LN2=0.07U WN2=0.7U
XI305 NET90 NET073 WLPCD2 S11000X8_SNAND LP2=0.07U WP2=0.42U LP1=0.07U WP1=0.42U LN1=0.07U
+WN1=0.21U LN2=0.07U WN2=0.21U
XI307 BLEQB WLPCD0 WLPCD4 S11000X8_SNAND LP2=0.07U WP2=1.75U LP1=0.07U WP1=3.5U LN1=0.07U
+WN1=4U LN2=0.07U WN2=4U
XI306 NET289 WLPCD1 BWEB_SU S11000X8_SNAND LP2=0.07U WP2=0.3U LP1=0.07U WP1=0.3U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI339 NET0219 DCLK WLPCD3 S11000X8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI186 NET163 NET93 NET073 S11000X8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI312 NET083 WLPCD0 S11000X8_SINV LP=0.10U WP=0.35U LN=0.10U WN=0.15U
XI73 GW_R GW_RB S11000X8_SINV LP=0.07U WP=1.4U LN=0.07U WN=0.7U
XI348 NET0100 GW_R S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI329 NET0153 WLPCD3 S11000X8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.15U
XI217 WLPCD1 WLPCD0 S11000X8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.28U
XI340 DLH NET0219 S11000X8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.7U
XI287 NET93 NET135 S11000X8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI327 NET141 NET139 S11000X8_SINV LP=0.18U WP=0.35U LN=0.18U WN=0.15U
XI286 NET135 PGB S11000X8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI134 SAE NET073 S11000X8_SINV LP=0.15U WP=0.7U LN=0.1U WN=0.35U
XI321 NET062 NET289 S11000X8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI264 WLPCD4 NET0153 S11000X8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI322 NET089 NET062 S11000X8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.2U
XI185 NET166 NET90 S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.28U
XI299 WLPCD2 NET100 S11000X8_SINV LP=0.07U WP=0.9U LN=0.07U WN=0.3U
XI298 NET100 WLPCD1 S11000X8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI207 NET_110 NET141 S11000X8_SINV LP=0.10U WP=0.7U LN=0.10U WN=0.28U
XI334 DLEQB NET095 S11000X8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
XI337 WLPCD3 WLPCD2 S11000X8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.25U
XI128 WLPCD0 NET085 S11000X8_SINV LP=0.07U WP=1.6U LN=0.07U WN=0.8U
XI315 NET085 WLP S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI333 NET095 BLEQB S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI311 NET088 NET083 S11000X8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
XI310 NET139 NET088 S11000X8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
**C50 WLPCD4 GND 2.8F
**C51 NET135 GND 0.45F
**C17 WLPCD1 GND 1.92F
**C33 NET139 GND 1F
**C15 NET0100 GND 0.57F
**C31 NET_110 GND 2.8F
**C13 NET073 GND 2.95F
**C10 NET095 GND 1.2F
**C11 NET0219 GND 1F
**C48 WLPCD2 GND 2.96F
**C47 NET166 GND 1F
**C26 BWEB_SU GND 1.6F
**C42 NET161 GND 2.1F
**C27 NET93 GND 1.6F
**C43 NET163 GND 0.85F
**C24 NET062 GND 0.7F
**C9 NET0153 GND 0.5F
**C8 WLPCD3 GND 1F
**C7 NET100 GND 0.55F
**C6 NET085 GND 0.6F
**C5 NET089 GND 2.4F
**C4 GW_R GND 4.29F
**C3 NET289 GND 1.1F
**C2 NET083 GND 0.5F
**C1 NET088 GND 1.1F
**C0 NET141 GND 0.7F
**C54 NET90 GND 0.45F
**C18 WLPCD0 GND 4F
.ENDS S11000X8_IO_RWCTRL_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IORWBLK_M16                                                          *
* LAST TIME SAVED: NOV 30 14:33:22 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IORWBLK_M16 BLEQB Q DL DLB AWTI BIST BWEB BWEBM D DCLK DM GW_RB WLP
XDIN AWTD BWEB_M NET46 BIST BWEB BWEBM D DM S11000X8_DIN
XSA Q AWTD AWTI DL DLB PGB PREB SAE S11000X8_SA
XIO_WRIN DL DLB NET46 DCLK_DATA NET041 WPG S11000X8_IO_WRIN_M16
XIO_RWCTRL BLEQB NET041 DCLK_DATA PGB PREB SAE WPG BWEB_M DCLK GW_RB WLP
+S11000X8_IO_RWCTRL_M16
**C3 WPG GND 5F
**C2 SAE GND 5F
**C8 NET041 GND 3.5F
**C4 PGB GND 5F
**C0 DCLK_DATA GND 2F
**C5 PREB GND 5F
**C6 BWEB_M GND 1.7F
**C7 AWTD GND 1.7F
**C1 NET46 GND 1.7F
.ENDS S11000X8_IORWBLK_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YSELX4                                                               *
* LAST TIME SAVED: DEC 12 10:42:39 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_YSELX4 YSEL[3] YSEL[2] YSEL[1] YSEL[0] Y10[3] Y10[2] Y10[1] Y10[0] Y432
**C76 NET15 GND 1.1F
**C77 NET26 GND 1.1F
**C79 NET43 GND 1.1F
**C81 NET40 GND 1.1F
XI73 YSEL[2] NET43 S11000X8_SINV LP=0.07U WP=0.84U LN=0.07U WN=0.41U
XI72 YSEL[1] NET26 S11000X8_SINV LP=0.07U WP=0.84U LN=0.07U WN=0.41U
XI61 YSEL[0] NET15 S11000X8_SINV LP=0.07U WP=0.84U LN=0.07U WN=0.41U
XI74 YSEL[3] NET40 S11000X8_SINV LP=0.07U WP=0.84U LN=0.07U WN=0.41U
MN4 NET40 Y10[3] NET12 GND NCH W=0.32U L=0.07U
MN1 NET15 Y10[0] NET12 GND NCH W=0.32U L=0.07U
MN3 NET43 Y10[2] NET12 GND NCH W=0.32U L=0.07U
MN0 NET12 Y432 GND GND NCH W=0.32U L=0.07U
MN2 NET26 Y10[1] NET12 GND NCH W=0.32U L=0.07U
MP6 VDD Y10[3] NET40 VDD PCH W=0.32U L=0.07U
MP7 VDD Y432 NET40 VDD PCH W=0.32U L=0.07U
MP5 VDD Y432 NET43 VDD PCH W=0.32U L=0.07U
MP3 VDD Y432 NET26 VDD PCH W=0.32U L=0.07U
MP4 VDD Y10[2] NET43 VDD PCH W=0.32U L=0.07U
MP1 VDD Y432 NET15 VDD PCH W=0.32U L=0.07U
MP2 VDD Y10[1] NET26 VDD PCH W=0.32U L=0.07U
MP0 VDD Y10[0] NET15 VDD PCH W=0.32U L=0.07U
.ENDS S11000X8_YSELX4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_M16                                                               *
* LAST TIME SAVED: NOV 10 11:38:59 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IO_M16 Q BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BL[8]
+BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[0] BLB[1] BLB[2] BLB[3]
+BLB[4] BLB[5] BLB[6] BLB[7] BLB[8] BLB[9] BLB[10] BLB[11] BLB[12] BLB[13] BLB[14]
+BLB[15] AWTI BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP Y10[3] Y10[2] Y10[1]
+Y10[0] Y32[3] Y32[2] Y32[1] Y32[0]
XIYPASS_15 BL[15] BLB[15] NET25 NET24 NET23 YSEL[15] S11000X8_IOYPASS_M16
XIYPASS_14 BL[14] BLB[14] NET25 NET24 NET23 YSEL[14] S11000X8_IOYPASS_M16
XIYPASS_13 BL[13] BLB[13] NET25 NET24 NET23 YSEL[13] S11000X8_IOYPASS_M16
XIYPASS_12 BL[12] BLB[12] NET25 NET24 NET23 YSEL[12] S11000X8_IOYPASS_M16
XIYPASS_11 BL[11] BLB[11] NET25 NET24 NET23 YSEL[11] S11000X8_IOYPASS_M16
XIYPASS_10 BL[10] BLB[10] NET25 NET24 NET23 YSEL[10] S11000X8_IOYPASS_M16
XIYPASS_9 BL[9] BLB[9] NET25 NET24 NET23 YSEL[9] S11000X8_IOYPASS_M16
XIYPASS_8 BL[8] BLB[8] NET25 NET24 NET23 YSEL[8] S11000X8_IOYPASS_M16
XIYPASS_7 BL[7] BLB[7] NET25 NET24 NET23 YSEL[7] S11000X8_IOYPASS_M16
XIYPASS_6 BL[6] BLB[6] NET25 NET24 NET23 YSEL[6] S11000X8_IOYPASS_M16
XIYPASS_5 BL[5] BLB[5] NET25 NET24 NET23 YSEL[5] S11000X8_IOYPASS_M16
XIYPASS_4 BL[4] BLB[4] NET25 NET24 NET23 YSEL[4] S11000X8_IOYPASS_M16
XIYPASS_3 BL[3] BLB[3] NET25 NET24 NET23 YSEL[3] S11000X8_IOYPASS_M16
XIYPASS_2 BL[2] BLB[2] NET25 NET24 NET23 YSEL[2] S11000X8_IOYPASS_M16
XIYPASS_1 BL[1] BLB[1] NET25 NET24 NET23 YSEL[1] S11000X8_IOYPASS_M16
XIYPASS_0 BL[0] BLB[0] NET25 NET24 NET23 YSEL[0] S11000X8_IOYPASS_M16
XI2 NET23 Q NET25 NET24 AWTI BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP
+S11000X8_IORWBLK_M16
XYSELX4_3 YSEL[15] YSEL[14] YSEL[13] YSEL[12] Y10[3] Y10[2] Y10[1] Y10[0]
+Y32[3] S11000X8_YSELX4
XYSELX4_2 YSEL[11] YSEL[10] YSEL[9] YSEL[8] Y10[3] Y10[2] Y10[1] Y10[0] Y32[2]
+S11000X8_YSELX4
XYSELX4_1 YSEL[7] YSEL[6] YSEL[5] YSEL[4] Y10[3] Y10[2] Y10[1] Y10[0] Y32[1]
+S11000X8_YSELX4
XYSELX4_0 YSEL[3] YSEL[2] YSEL[1] YSEL[0] Y10[3] Y10[2] Y10[1] Y10[0] Y32[0]
+S11000X8_YSELX4
.ENDS S11000X8_IO_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_WRIN_M8                                                           *
* LAST TIME SAVED: SEP 28 10:50:28 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IO_WRIN_M8 DL DLB D DCLK DLEQB WPG
XLH_DCLK_M8 D1B DCLK D S11000X8_LH_DCLK
MP7 DL DLEQB VDD VDD PCH W=1U L=0.07U
MP8 VDD DLEQB DLB VDD PCH W=1U L=0.07U
MN2 VDD D1 D2B VDD PCH W=2.5U L=0.07U
MN0 VDD D1B D2 VDD PCH W=2.5U L=0.07U
MN5 DLB WPG D2B GND NCH W=2.5U L=0.07U
MN4 D2 WPG DL GND NCH W=2.5U L=0.07U
MN3 D2B D1 GND GND NCH W=5U L=0.07U
MN1 D2 D1B GND GND NCH W=5U L=0.07U
XI69 D1 D1B S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
**C11 D1B GND 4.2F
**C6 D1 GND 2.6F
**C7 D2B GND 4.5F
**C8 D2 GND 4.5F
.ENDS S11000X8_IO_WRIN_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_RWCTRL_M8                                                         *
* LAST TIME SAVED: OCT  6 16:44:21 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IO_RWCTRL_M8 BLEQB DLEQB DLH PGB PREB SAE WPG BWEB DCLK GW_RB WLP
X_LH_BWEB BWEB_SU DLH BWEB S11000X8_LH_BWEB
XI289 PREB NET0100 NET161 S11000X8_SNOR LP1=0.07U WP1=1.2U LP2=0.07U WP2=1.2U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI288 NET161 WLPCD2 NET163 S11000X8_SNOR LP1=0.07U WP1=0.35U LP2=0.07U WP2=0.35U LN2=0.07U
+WN2=0.3U LN1=0.07U WN1=0.3U
XI249 WPG GW_R NET089 S11000X8_SNOR LP1=0.07U WP1=1.0U LP2=0.07U WP2=1.0U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI133 NET073 WLPCD0 NET_110 GW_R S11000X8_SNAND3 LP3=0.07U WP3=1.75U LP2=0.07U WP2=1.75U
+LP1=0.07U WP1=1.75U LN1=0.07U WN1=1.2U LN2=0.07U WN2=1.2U LN3=0.07U WN3=1.2U
XI250 PGB NET166 GW_R S11000X8_SNAND LP2=0.07U WP2=0.84U LP1=0.07U WP1=0.84U LN1=0.07U
+WN1=0.7U LN2=0.07U WN2=0.7U
XI305 NET90 NET073 WLPCD2 S11000X8_SNAND LP2=0.07U WP2=0.42U LP1=0.07U WP1=0.42U LN1=0.07U
+WN1=0.21U LN2=0.07U WN2=0.21U
XI307 BLEQB WLPCD0 WLPCD4 S11000X8_SNAND LP2=0.07U WP2=1.75U LP1=0.07U WP1=3.5U LN1=0.07U
+WN1=4U LN2=0.07U WN2=4U
XI306 NET289 WLPCD1 BWEB_SU S11000X8_SNAND LP2=0.07U WP2=0.3U LP1=0.07U WP1=0.3U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI339 NET0219 DCLK WLPCD3 S11000X8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI186 NET163 NET93 NET073 S11000X8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI312 NET083 WLPCD0 S11000X8_SINV LP=0.10U WP=0.35U LN=0.10U WN=0.15U
XI73 GW_R GW_RB S11000X8_SINV LP=0.07U WP=1.4U LN=0.07U WN=0.7U
XI348 NET0100 GW_R S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI329 NET0153 WLPCD3 S11000X8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.15U
XI217 WLPCD1 WLPCD0 S11000X8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.28U
XI340 DLH NET0219 S11000X8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.7U
XI287 NET93 NET135 S11000X8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI327 NET141 NET139 S11000X8_SINV LP=0.18U WP=0.35U LN=0.18U WN=0.15U
XI286 NET135 PGB S11000X8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI134 SAE NET073 S11000X8_SINV LP=0.15U WP=0.7U LN=0.1U WN=0.35U
XI321 NET062 NET289 S11000X8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI264 WLPCD4 NET0153 S11000X8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI322 NET089 NET062 S11000X8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.2U
XI185 NET166 NET90 S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.28U
XI299 WLPCD2 NET100 S11000X8_SINV LP=0.07U WP=0.9U LN=0.07U WN=0.3U
XI298 NET100 WLPCD1 S11000X8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI207 NET_110 NET141 S11000X8_SINV LP=0.10U WP=0.7U LN=0.10U WN=0.28U
XI334 DLEQB NET095 S11000X8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
XI337 WLPCD3 WLPCD2 S11000X8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.25U
XI128 WLPCD0 NET085 S11000X8_SINV LP=0.07U WP=1.6U LN=0.07U WN=0.8U
XI315 NET085 WLP S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI333 NET095 BLEQB S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI311 NET088 NET083 S11000X8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
XI310 NET139 NET088 S11000X8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
**C50 WLPCD4 GND 2.8F
**C51 NET135 GND 0.45F
**C17 WLPCD1 GND 1.92F
**C33 NET139 GND 1F
**C15 NET0100 GND 0.57F
**C31 NET_110 GND 2.8F
**C13 NET073 GND 2.95F
**C10 NET095 GND 1.2F
**C11 NET0219 GND 1F
**C48 WLPCD2 GND 2.96F
**C47 NET166 GND 1F
**C26 BWEB_SU GND 1.6F
**C42 NET161 GND 2.1F
**C27 NET93 GND 1.6F
**C43 NET163 GND 0.85F
**C24 NET062 GND 0.7F
**C9 NET0153 GND 0.5F
**C8 WLPCD3 GND 1F
**C7 NET100 GND 0.55F
**C6 NET085 GND 0.6F
**C5 NET089 GND 2.4F
**C4 GW_R GND 4.29F
**C3 NET289 GND 1.1F
**C2 NET083 GND 0.5F
**C1 NET088 GND 1.1F
**C0 NET141 GND 0.7F
**C54 NET90 GND 0.45F
**C18 WLPCD0 GND 4F
.ENDS S11000X8_IO_RWCTRL_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IORWBLK_M8                                                           *
* LAST TIME SAVED: DEC 14 17:21:00 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IORWBLK_M8 BLEQB Q DL DLB AWTI BIST BWEB BWEBM D DCLK DM GW_RB WLP
XDIN AWTD BWEB_M NET42 BIST BWEB BWEBM D DM S11000X8_DIN
XSA Q AWTD AWTI DL DLB PGB PREB SAE S11000X8_SA
XIO_WRIN DL DLB NET42 DCLK_DATA NET041 WPG S11000X8_IO_WRIN_M8
XIO_RWCTRL BLEQB NET041 DCLK_DATA PGB PREB SAE WPG BWEB_M DCLK GW_RB WLP
+S11000X8_IO_RWCTRL_M8
**C3 WPG GND 1.7F
**C2 SAE GND 3F
**C8 NET041 GND 1.5F
**C4 PGB GND 4.3F
**C0 DCLK_DATA GND 4.7F
**C5 PREB GND 2.1F
**C7 AWTD GND 1.7F
**C6 BWEB_M GND 1.7F
**C1 NET42 GND 1.7F
.ENDS S11000X8_IORWBLK_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IOYPASS_M8                                                           *
* LAST TIME SAVED: DEC 14 17:22:46 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IOYPASS_M8 BL BLB DL DLB BLEQB YSEL
**C19 NET47 GND 0.97F
*MN0 BL YSEL DL GND NCH W=0.8U L=0.06U
MN0 BL YSEL DL GND NCH W=0.89U L=0.06U
*MN1 BLB YSEL DLB GND NCH W=0.8U L=0.06U
MN1 BLB YSEL DLB GND NCH W=0.89U L=0.06U
MP2 BLB BLEQB BL VDD PCH W=2U L=0.06U
MP0 BL NET47 DL VDD PCH W=0.8U L=0.06U
MP3 VDD BLEQB BLB VDD PCH W=2U L=0.06U
MP1 BLB NET47 DLB VDD PCH W=0.8U L=0.06U
MP4 BL BLEQB VDD VDD PCH W=2U L=0.06U
XI9 NET47 YSEL S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.24U
.ENDS S11000X8_IOYPASS_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_M8                                                                *
* LAST TIME SAVED: DEC  2 19:25:13 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IO_M8 Q BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] BLB[1]
+BLB[2] BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] AWTI BIST_BUF BWEB BWEBM D DCLK DM
+GW_RB WLP Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0]
**CI6_7 YSEL[7] GND 1.7F
**CI6_6 YSEL[6] GND 1.7F
**CI6_5 YSEL[5] GND 1.7F
**CI6_4 YSEL[4] GND 1.7F
**CI6_3 YSEL[3] GND 1.7F
**CI6_2 YSEL[2] GND 1.7F
**CI6_1 YSEL[1] GND 1.7F
**CI6_0 YSEL[0] GND 1.7F
**CI7 NET31 GND 13F
**CI9 NET32 GND 8.13F
**CI11 NET33 GND 8.09F
XI2 NET31 Q NET33 NET32 AWTI BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP S11000X8_IORWBLK_M8
XYSELX4_1 YSEL[7] YSEL[6] YSEL[5] YSEL[4] Y10[3] Y10[2] Y10[1] Y10[0] Y32[1]
+S11000X8_YSELX4
XYSELX4_0 YSEL[3] YSEL[2] YSEL[1] YSEL[0] Y10[3] Y10[2] Y10[1] Y10[0] Y32[0]
+S11000X8_YSELX4
XIYPASS_7 BL[7] BLB[7] NET33 NET32 NET31 YSEL[7] S11000X8_IOYPASS_M8
XIYPASS_6 BL[6] BLB[6] NET33 NET32 NET31 YSEL[6] S11000X8_IOYPASS_M8
XIYPASS_5 BL[5] BLB[5] NET33 NET32 NET31 YSEL[5] S11000X8_IOYPASS_M8
XIYPASS_4 BL[4] BLB[4] NET33 NET32 NET31 YSEL[4] S11000X8_IOYPASS_M8
XIYPASS_3 BL[3] BLB[3] NET33 NET32 NET31 YSEL[3] S11000X8_IOYPASS_M8
XIYPASS_2 BL[2] BLB[2] NET33 NET32 NET31 YSEL[2] S11000X8_IOYPASS_M8
XIYPASS_1 BL[1] BLB[1] NET33 NET32 NET31 YSEL[1] S11000X8_IOYPASS_M8
XIYPASS_0 BL[0] BLB[0] NET33 NET32 NET31 YSEL[0] S11000X8_IOYPASS_M8
.ENDS S11000X8_IO_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_WRIN_M4                                                           *
* LAST TIME SAVED: DEC 14 16:50:06 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IO_WRIN_M4 DL DLB D DCLK DLEQB WPG
XLH_DCLK_M8 D1B DCLK D S11000X8_LH_DCLK
MP7 DL DLEQB VDD VDD PCH W=1U L=0.07U
MP8 VDD DLEQB DLB VDD PCH W=1U L=0.07U
MN2 VDD D1 D2B VDD PCH W=2.5U L=0.07U
MN0 VDD D1B D2 VDD PCH W=2.5U L=0.07U
MN5 DLB WPG D2B GND NCH W=2.5U L=0.07U
MN4 D2 WPG DL GND NCH W=2.5U L=0.07U
MN3 D2B D1 GND GND NCH W=5U L=0.07U
MN1 D2 D1B GND GND NCH W=5U L=0.07U
XI69 D1 D1B S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
**C11 D1B GND 5.983F
**C6 D1 GND 3.851F
**C7 D2B GND 2.669F
**C8 D2 GND 3.188F
.ENDS S11000X8_IO_WRIN_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_RWCTRL_M4                                                         *
* LAST TIME SAVED: DEC 14 16:50:07 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IO_RWCTRL_M4 BLEQB DLEQB DLH PGB PREB SAE WPG BWEB DCLK GW_RB WLP
X_LH_BWEB BWEB_SU DLH BWEB S11000X8_LH_BWEB
XI289 PREB NET0100 NET161 S11000X8_SNOR LP1=0.07U WP1=1.2U LP2=0.07U WP2=1.2U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI288 NET161 WLPCD2 NET163 S11000X8_SNOR LP1=0.07U WP1=0.35U LP2=0.07U WP2=0.35U LN2=0.07U
+WN2=0.3U LN1=0.07U WN1=0.3U
XI249 WPG GW_R NET089 S11000X8_SNOR LP1=0.07U WP1=1.0U LP2=0.07U WP2=1.0U LN2=0.07U
+WN2=0.4U LN1=0.07U WN1=0.4U
XI133 NET073 WLPCD0 NET_110 GW_R S11000X8_SNAND3 LP3=0.07U WP3=1.75U LP2=0.07U WP2=1.75U
+LP1=0.07U WP1=1.75U LN1=0.07U WN1=1.2U LN2=0.07U WN2=1.2U LN3=0.07U WN3=1.2U
XI250 PGB NET166 GW_R S11000X8_SNAND LP2=0.07U WP2=0.84U LP1=0.07U WP1=0.84U LN1=0.07U
+WN1=0.7U LN2=0.07U WN2=0.7U
XI305 NET90 NET073 WLPCD2 S11000X8_SNAND LP2=0.07U WP2=0.42U LP1=0.07U WP1=0.42U LN1=0.07U
+WN1=0.21U LN2=0.07U WN2=0.21U
XI307 BLEQB WLPCD0 WLPCD4 S11000X8_SNAND LP2=0.07U WP2=1.75U LP1=0.07U WP1=3.5U LN1=0.07U
+WN1=1U LN2=0.07U WN2=1U
XI306 NET289 WLPCD1 BWEB_SU S11000X8_SNAND LP2=0.07U WP2=0.3U LP1=0.07U WP1=0.3U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI339 NET0219 DCLK WLPCD3 S11000X8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI186 NET163 NET93 NET073 S11000X8_SNAND LP2=0.07U WP2=0.35U LP1=0.07U WP1=0.35U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI312 NET083 WLPCD0 S11000X8_SINV LP=0.10U WP=0.35U LN=0.10U WN=0.15U
XI73 GW_R GW_RB S11000X8_SINV LP=0.07U WP=1.4U LN=0.07U WN=0.7U
XI348 NET0100 GW_R S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI329 NET0153 WLPCD3 S11000X8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.15U
XI217 WLPCD1 WLPCD0 S11000X8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.28U
XI340 DLH NET0219 S11000X8_SINV LP=0.07U WP=0.7U LN=0.07U WN=0.7U
XI287 NET93 NET135 S11000X8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI327 NET141 NET139 S11000X8_SINV LP=0.18U WP=0.35U LN=0.18U WN=0.15U
XI286 NET135 PGB S11000X8_SINV LP=0.07U WP=0.15U LN=0.07U WN=0.15U
XI134 SAE NET073 S11000X8_SINV LP=0.15U WP=0.7U LN=0.1U WN=0.35U
XI321 NET062 NET289 S11000X8_SINV LP=0.07U WP=0.30U LN=0.07U WN=0.15U
XI264 WLPCD4 NET0153 S11000X8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI322 NET089 NET062 S11000X8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.2U
XI185 NET166 NET90 S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.28U
XI299 WLPCD2 NET100 S11000X8_SINV LP=0.07U WP=0.9U LN=0.07U WN=0.3U
XI298 NET100 WLPCD1 S11000X8_SINV LP=0.07U WP=0.35U LN=0.07U WN=0.35U
XI207 NET_110 NET141 S11000X8_SINV LP=0.10U WP=0.7U LN=0.10U WN=0.28U
XI334 DLEQB NET095 S11000X8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
XI337 WLPCD3 WLPCD2 S11000X8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.25U
XI128 WLPCD0 NET085 S11000X8_SINV LP=0.07U WP=1.6U LN=0.07U WN=0.8U
XI315 NET085 WLP S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI333 NET095 BLEQB S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI311 NET088 NET083 S11000X8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
XI310 NET139 NET088 S11000X8_SINV LP=0.35U WP=0.35U LN=0.35U WN=0.15U
**C50 WLPCD4 GND 1.317F
**C51 NET135 GND 0.555F
**C17 WLPCD1 GND 1.524F
**C33 NET139 GND 0.850F
**C15 NET0100 GND 2.197F
**C31 NET_110 GND 2.187F
**C13 NET073 GND 3.990F
**C10 NET095 GND 0.690F
**C11 NET0219 GND 1.025F
**C48 WLPCD2 GND 3.190F
**C47 NET166 GND 0.853F
**C26 BWEB_SU GND 2.568F
**C42 NET161 GND 0.935F
**C27 NET93 GND 0.533F
**C43 NET163 GND 1.781F
**C24 NET062 GND 0.737F
**C9 NET0153 GND 1.066F
**C8 WLPCD3 GND 3.831F
**C7 NET100 GND 0.733F
**C6 NET085 GND 1.719F
**C5 NET089 GND 0.959F
**C4 GW_R GND 6.770F
**C3 NET289 GND 0.760F
**C2 NET083 GND 0.902F
**C1 NET088 GND 0.616F
**C0 NET141 GND 0.837F
**C54 NET90 GND 2.157F
**C18 WLPCD0 GND 7.540F
.ENDS S11000X8_IO_RWCTRL_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IORWBLK_M4                                                           *
* LAST TIME SAVED: DEC  8 17:33:56 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IORWBLK_M4 BLEQB Q DL DLB AWTI BIST BWEB BWEBM D DCLK DM GW_RB WLP
XDIN AWTD BWEB_M NET47 BIST BWEB BWEBM D DM S11000X8_DIN
XIO_WRIN DL DLB NET47 DCLK_DATA NET041 WPG S11000X8_IO_WRIN_M4
XIO_RWCTRL BLEQB NET041 DCLK_DATA PGB PREB SAE WPG BWEB_M DCLK GW_RB WLP
+S11000X8_IO_RWCTRL_M4
XSA Q AWTD AWTI DL DLB PGB PREB SAE S11000X8_SA
**C3 WPG GND 3.447F
**C2 SAE GND 5.928F
**C9 BLEQB GND 4.8F
**C8 NET041 GND 1.500F
**C4 PGB GND 6.882F
**C0 DCLK_DATA GND 6.355F
**C5 PREB GND 5.536F
**C6 BWEB_M GND 1.497F
**C7 AWTD GND 6.791F
**C1 NET47 GND 5.644F
.ENDS S11000X8_IORWBLK_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IOYPASS_M4                                                           *
* LAST TIME SAVED: DEC 14 16:50:08 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IOYPASS_M4 BL BLB DL DLB BLEQB YSEL
**C1 NET47 GND 1.979F
*MN0 BL YSEL DL GND NCH W=0.8U L=0.06U
MN0 BL YSEL DL GND NCH W=0.89U L=0.06U
*MN1 BLB YSEL DLB GND NCH W=0.8U L=0.06U
MN1 BLB YSEL DLB GND NCH W=0.89U L=0.06U
MP2 BLB BLEQB BL VDD PCH W=2U L=0.06U
MP0 BL NET47 DL VDD PCH W=0.8U L=0.06U
MP3 VDD BLEQB BLB VDD PCH W=2U L=0.06U
MP1 BLB NET47 DLB VDD PCH W=0.8U L=0.06U
MP4 BL BLEQB VDD VDD PCH W=2U L=0.06U
XI9 NET47 YSEL S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.24U
.ENDS S11000X8_IOYPASS_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: IO_M4                                                                *
* LAST TIME SAVED: DEC 15 14:54:17 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_IO_M4 Q BL[0] BL[1] BL[2] BL[3] BLB[0] BLB[1] BLB[2] BLB[3] AWTI
+BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP Y10[3] Y10[2] Y10[1] Y10[0]
XI2 NET23 Q NET25 NET24 AWTI BIST_BUF BWEB BWEBM D DCLK DM GW_RB WLP S11000X8_IORWBLK_M4
XIYPASS_3 BL[3] BLB[3] NET25 NET24 NET23 Y10[3] S11000X8_IOYPASS_M4
XIYPASS_2 BL[2] BLB[2] NET25 NET24 NET23 Y10[2] S11000X8_IOYPASS_M4
XIYPASS_1 BL[1] BLB[1] NET25 NET24 NET23 Y10[1] S11000X8_IOYPASS_M4
XIYPASS_0 BL[0] BLB[0] NET25 NET24 NET23 Y10[0] S11000X8_IOYPASS_M4
**C4 NET23 GND 15.052F
**C1 NET25 GND 9.518F
**C0 NET24 GND 9.433F
.ENDS S11000X8_IO_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SINV_HVT                                                             *
* LAST TIME SAVED: SEP 21 15:49:08 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_SINV_HVT Y A LP=0.06U WP=0.3U LN=0.06U WN=0.15U
M0 Y A GND GND NCH_HVT W=WN L=LN
M1 VDD A Y VDD PCH_HVT W=WP L=LP
.ENDS S11000X8_SINV_HVT


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V3                                                             *
* LAST TIME SAVED: DEC 14 16:49:42 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_DELAY_V3 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET28 TSEL IN S11000X8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI163 OUT_B NET28 S11000X8_SINV_HVT LP=0.32U WP=0.6U LN=0.32U WN=0.3U
**C153 NET28 GND 0.7F
.ENDS S11000X8_DELAY_V3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V2                                                             *
* LAST TIME SAVED: DEC 14 16:49:31 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_DELAY_V2 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET44 TSEL IN S11000X8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI165 OUT_B NET44 S11000X8_SINV_HVT LP=0.18U WP=0.6U LN=0.18U WN=0.3U
**C153 NET44 GND 0.7F
.ENDS S11000X8_DELAY_V2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V1                                                             *
* LAST TIME SAVED: DEC 14 16:49:18 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_DELAY_V1 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET27 TSEL IN S11000X8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI141 OUT_B NET27 S11000X8_SINV_HVT LP=0.12U WP=0.6U LN=0.12U WN=0.3U
**C151 NET27 GND 1.1F
.ENDS S11000X8_DELAY_V1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_CEB                                                               *
* LAST TIME SAVED: DEC 14 16:50:09 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_LH_CEB Q CP D
XI26 D P2 CP INCP S11000X8_TRANSGATE LP=0.07U WP=1U LN=0.07U WN=1U
MN12 GND Q NET39 GND NCH W=0.15U L=0.07U
MN11 NET39 INCP P2 GND NCH W=0.15U L=0.07U
MP4 NET69 Q VDD VDD PCH W=0.28U L=0.07U
MP5 P2 CP NET69 VDD PCH W=0.28U L=0.07U
XI33 Q P2 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI29 INCP CP S11000X8_SINV LP=0.07U WP=0.6U LN=0.07U WN=0.3U
**C1 P2 GND 1.955F
**C0 INCP GND 0.828F
.ENDS S11000X8_LH_CEB


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: PREBUF                                                               *
* LAST TIME SAVED: DEC 14 16:50:09 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_PREBUF SCLK_X SCLK_Y CEB CLK WLPX
X_LH_CEB H1 CK2 NET0309 S11000X8_LH_CEB
XI345 CK2 NET0179 H1 H0 S11000X8_TRANSGATE LP=0.06U WP=3.5U LN=0.06U WN=3.5U
MP4 NET0179 H1 VDD VDD PCH W=2U L=0.06U
XI358 CK2 NET0130 CLK S11000X8_SNOR LP1=0.06U WP1=3U LP2=0.06U WP2=3U LN2=0.06U WN2=3U
+LN1=0.06U WN1=3U
XI356 SCLK_Y NET0179 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=5U M=1
XI382 SCLK_X NET0179 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=5U M=2
XI353 H0 H1 S11000X8_SINV LP=0.06U WP=1U LN=0.06U WN=0.5U
XI354 NET0309 NET0297 S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI357 NET0302 NET0304 S11000X8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI359 NET0304 WLPX S11000X8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI361 NET0130 NET0302 S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI404 NET0297 CEB S11000X8_SINV LP=0.10U WP=0.3U LN=0.10U WN=0.15U
**C8 NET0179 GND 15.756F
**C9 H1 GND 5.364F
**C10 NET0309 GND 1.493F
**C12 H0 GND 1.999F
**C14 NET0297 GND 0.677F
**C39 NET0130 GND 2.062F
**C37 NET0304 GND 0.598F
**C38 NET0302 GND 0.748F
**C43 CK2 GND 7.480F
.ENDS S11000X8_PREBUF


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DFFQ_WEB                                                             *
* LAST TIME SAVED: DEC 14 16:50:10 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_DFFQ_WEB Q CP D
XI30 INV2 P2 INCP CP S11000X8_TRANSGATE LP=0.07U WP=2U LN=0.07U WN=1U
MN17 NET38 Q GND GND NCH W=0.3U L=0.07U
MN15 NET44 INV2 GND GND NCH W=0.2U L=0.07U
MN16 P2 CP NET38 GND NCH W=0.3U L=0.07U
MN14 INV1 INCP NET44 GND NCH W=0.2U L=0.07U
MN13 NET54 D GND GND NCH W=0.3U L=0.07U
MN7 INV1 CP NET54 GND NCH W=0.3U L=0.07U
MP10 NET68 INCP P2 VDD PCH W=0.6U L=0.07U
MP0 VDD D NET78 VDD PCH W=0.6U L=0.07U
MP7 VDD INV2 NET74 VDD PCH W=0.4U L=0.07U
MP6 NET78 INCP INV1 VDD PCH W=0.6U L=0.07U
MP8 NET74 CP INV1 VDD PCH W=0.4U L=0.07U
MP9 VDD Q NET68 VDD PCH W=0.6U L=0.07U
XI31 Q P2 S11000X8_SINV LP=0.07U WP=10U LN=0.07U WN=5U
XI33 INCP CP S11000X8_SINV LP=0.07U WP=1.00U LN=0.07U WN=0.35U
XI29 INV2 INV1 S11000X8_SINV LP=0.07U WP=3.0U LN=0.07U WN=1.5U
**C0 INV1 GND 2.338F
**C1 INCP GND 2.995F
**C2 INV2 GND 2.715F
**C3 P2 GND 5.625F
.ENDS S11000X8_DFFQ_WEB


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CLKBUF                                                               *
* LAST TIME MODIFIED: JULY 24 09:50:10 2006                                       *
*******************************************************************************
.SUBCKT S11000X8_CLKBUF DCLK GW_RB CEB CLK WEB
X_LH_DCLK H3 CK_WEB NET111 S11000X8_LH_DCLK
X_DFFQ_WEB NET69 CK_WEB SH S11000X8_DFFQ_WEB
***------------REMOVE------------------------------------------------------****
**XI273 CLK NET94 H3 H2 TRANSGATE LP=0.06U WP=2.1U LN=0.06U WN=2.1U
**MN10 NET94 H2 GND GND NCH W=0.2U L=0.1U
***------------ADD BELOW MOS------------------------------------------------------****
MP10 DCLK0 H3 VDD VDD PCH W=0.4U L=0.06U
XI1274 NET94 DCLK0 S11000X8_SINV LP=0.06U WP=4U LN=0.06U WN=2U 
MP1 VDD CLK NET001 VDD PCH W=1U L=0.06U
MP2 NET001 H2 DCLK0 VDD PCH W=1U L=0.06U
MN1 NET002 H3 DCLK0 GND NCH W=1U L=0.06U
MN2 GND CLK NET002 GND NCH W=1U L=0.06U
***-----------------------------------------------------------------------------*********
XI271 SH CEB WEB S11000X8_SNOR LP1=0.07U WP1=0.45U LP2=0.07U WP2=0.45U LN2=0.07U WN2=0.15U
+LN1=0.07U WN1=0.15U
XI246 GW_RB NET69 S11000X8_SINV LP=0.06U WP=9U LN=0.06U WN=4.5U M=2
XI280 H2 H3 S11000X8_SINV LP=0.06U WP=0.35U LN=0.06U WN=0.15U
XI277 NET111 SH S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI202 CK_WEB CLK S11000X8_SINV LP=0.06U WP=0.8U LN=0.06U WN=0.8U
XI274 DCLK NET94 S11000X8_SINV LP=0.06U WP=8U LN=0.06U WN=8U M=2
**C43 SH GND 4.641F
**C18 CK_WEB GND 7.391F
**C19 NET69 GND 12.723F
**C21 NET94 GND 13.840F
**C24 H3 GND 4.176F
**C26 NET111 GND 1.130F
**C27 SH GND 4.641F
**C25 H2 GND 1.913F
.ENDS S11000X8_CLKBUF


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M16V1                                                         *
* LAST TIME SAVED: DEC  1 14:30:39 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_WLPGEN_M16V1 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK
+TM TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 NET122 D02 SEL[3] SELN[3] SELN[2] S11000X8_DELAY_V3
XI337 D02 NET122 D01 SEL[2] SELN[2] SELN[1] S11000X8_DELAY_V2
XI326 D01 NET122 NET0214 SEL[1] SELN[1] SELN[0] S11000X8_DELAY_V1
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S11000X8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S11000X8_CLKBUF
**XI324 NET122 NET0214 SEL[0] SELN[0] TRANSGATE LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI324 NET122 NET1227 SEL[0] SELN[0] S11000X8_TRANSGATE LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI238 D1 T0 NET132 CLK_K S11000X8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S11000X8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET169 CLK_KB CLK S11000X8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN7 NET96 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET097 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET096 GND NCH W=5U L=0.06U
MN0 NET096 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET96 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET0198 NET097 GND NCH W=5U L=0.07U
MP5 VDD TME NET0108 VDD PCH W=10U L=0.06U M=2
MP9 NET80 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET0119 NET0198 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET0108 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET80 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET0119 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI219 NET169 WLP_RESET WLPSTART S11000X8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI482 WLP_RESET NET122 NET210 S11000X8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U LN1=0.06U
+WN1=1.0U LN2=0.06U WN2=1.0U
XI328 SELN[0] SEL0N SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S11000X8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI383 NET0198 WLPTEST S11000X8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI386 TRWLPB TRWLP S11000X8_SINV LP=0.2U WP=1.0U LN=0.2U WN=0.4U
XI471 SEL[3] SELN[3] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET0323 S11000X8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET0321 CEB S11000X8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET0348 WLPSTART S11000X8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET0354 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET0354 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI371 NET0323 NET0321 S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI292 NET0214 TRWLPB S11000X8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI283 CLK_KB CLK S11000X8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
**XI493 NET209 NET122 SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI493 NET1227 NET0214 S11000X8_SINV LP=0.06U WP=0.755U LN=0.06U WN=0.2U
XI495 NET213 NET208 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI296 CLK_K NET132 S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI297 NET132 CLK S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**XI494 NET208 NET209 SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI494 NET208 NET122 S11000X8_SINV LP=0.06U WP=0.755U LN=0.06U WN=0.2U
XI473 SEL1 SEL1N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI497 NET210 TRWLP S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI315 TME TMEB S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI496 NET211 NET213 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
**CI414 D03 GND 0.7F
**C36 TRWLPB GND 5.4F
**CI428 D02 GND 1.2F
**C40 NET0354 GND 5.6F
**CI410 SEL0 GND 2.1F
**CI446 TME GND 5.5F
**CI426 D01 GND 1.3F
**CI420 SEL0N GND 2.9F
**CI434 NET0214 GND 1.5F
**CI448 TMEB GND 6.1F
**C0 T2 GND 6.1F
**C4 NET132 GND 0.7F
**CI418 SEL1 GND 2.7F
**C34 WLPSTART GND 13.1F
**C35 NET0348 GND 8.2F
**CI432 NET0198 GND 5.2F
**C30 NET0323 GND 0.7F
**C15 NET0321 GND 0.7F
**CI422 SEL1N GND 2.8F
**C32 D1 GND 1.4F
**C1 T1 GND 3.2F
**C5 CLK_K GND 0.8F
**CI444 SELN[0] GND 3.9F
**C22 CLK_KB GND 2.2F
**CI442 SEL[0] GND 4.1F
**C33 T0 GND 1.0F
**C31 NET169 GND 5.6F
**C2 WLP_RESET GND 5.5F
.ENDS S11000X8_WLPGEN_M16V1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CEBBISMX                                                             *
* LAST TIME SAVED: NOV 30 14:35:28 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_CEBBISMX MXOUT A AM BISTC BISTT
**C0 GND NET30 1.033F
XI5 MXOUT NET30 S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
MP15 Z21 BISTT NET30 VDD PCH W=0.5U L=0.06U
MP14 VDD A Z21 VDD PCH W=0.5U L=0.06U
MP7 VDD AM Z22 VDD PCH W=0.5U L=0.06U
MP6 Z22 BISTC NET30 VDD PCH W=0.5U L=0.06U
MN15 NET30 BISTC Z23 GND NCH W=0.25U L=0.06U
MN14 NET30 BISTT Z24 GND NCH W=0.25U L=0.06U
MN13 Z23 A GND GND NCH W=0.25U L=0.06U
MN6 Z24 AM GND GND NCH W=0.25U L=0.06U
.ENDS S11000X8_CEBBISMX


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AWTD_M16                                                             *
* LAST TIME SAVED: OCT  4 16:21:02 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_AWTD_M16 AWTI AWT
XINV0 AWTI Z1 S11000X8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI9 Z1 AWT S11000X8_SINV LP=0.07U WP=3U LN=0.07U WN=1.5U
.ENDS S11000X8_AWTD_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISTD_M16                                                            *
* LAST TIME SAVED: OCT  4 16:22:00 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BISTD_M16 BISTC BISTT BIST
XI13 BISTT BISTC S11000X8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI14 BISTC BIST S11000X8_SINV LP=0.07U WP=3.2U LN=0.07U WN=1.6U
.ENDS S11000X8_BISTD_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISIN_M16                                                            *
* LAST TIME SAVED: DEC  1 14:16:28 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BISIN_M16 AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM
XCEBMX CEBX CEB CEBM BISTC BIST_BUF S11000X8_CEBBISMX
XWEBMX WEBX WEB WEBM BISTC BIST_BUF S11000X8_CEBBISMX
XAWTD AWTI AWT S11000X8_AWTD_M16
XBISTD BISTC BIST_BUF BIST S11000X8_BISTD_M16
.ENDS S11000X8_BISIN_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: SRAM_TIEL                                                            *
* LAST TIME SAVED: MAY 16 14:03:38 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_SRAM_TIEL Z
XI49 Z NET14 S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=4U
MN1 GND NET14 NET32 GND NCH W=0.15U L=0.07U
MN0 NET32 NET32 GND GND NCH W=0.15U L=0.07U
MP0 VDD NET32 NET14 VDD PCH W=0.3U L=0.07U
.ENDS S11000X8_SRAM_TIEL


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_YPD_M16                                                           *
* LAST TIME SAVED: SEP 30 15:10:52 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_LH_YPD_M16 Q CP D
XI26 D P2 INCPN CP S11000X8_TRANSGATE LP=0.07U WP=2U LN=0.07U WN=2U
MN0 GND Q NET38 GND NCH W=0.2U L=0.07U
MN1 NET38 CP P2 GND NCH W=0.2U L=0.07U
MP4 NET49 Q VDD VDD PCH W=0.5U L=0.07U
MP5 P2 INCPN NET49 VDD PCH W=0.5U L=0.07U
XI23 Q P2 S11000X8_SINV LP=0.07U WP=8U LN=0.07U WN=4U
XI29 INCPN CP S11000X8_SINV LP=0.07U WP=1.2U LN=0.07U WN=0.6U
**C2 P2 GND 3F
**C3 INCPN GND 1.5F
.ENDS S11000X8_LH_YPD_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPRE10_M16                                                           *
* LAST TIME SAVED: DEC 13 14:07:14 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_YPRE10_M16 Y10[3] Y10[2] Y10[1] Y10[0] BISTT SCLK Y[1] Y[0] YM[1] YM[0]
MP0 NET43 BISTC Y1N VDD PCH W=0.3U L=0.07U
MP15 NET40 BISTT Y0N VDD PCH W=0.3U L=0.07U
MP14 VDD Y[0] NET40 VDD PCH W=0.3U L=0.07U
MP7 VDD YM[0] NET31 VDD PCH W=0.3U L=0.07U
MP6 NET31 BISTC Y0N VDD PCH W=0.3U L=0.07U
MP1 VDD YM[1] NET43 VDD PCH W=0.3U L=0.07U
MP2 VDD Y[1] NET22 VDD PCH W=0.3U L=0.07U
MP3 NET22 BISTT Y1N VDD PCH W=0.3U L=0.07U
MN3 Y1N BISTC NET46 GND NCH W=0.15U L=0.07U
MN2 Y1N BISTT NET49 GND NCH W=0.15U L=0.07U
MN15 Y0N BISTC NET55 GND NCH W=0.15U L=0.07U
MN14 Y0N BISTT NET52 GND NCH W=0.15U L=0.07U
MN13 NET55 Y[0] GND GND NCH W=0.15U L=0.07U
MN6 NET52 YM[0] GND GND NCH W=0.15U L=0.07U
MN0 NET49 YM[1] GND GND NCH W=0.15U L=0.07U
MN1 NET46 Y[1] GND GND NCH W=0.15U L=0.07U
XLH_YPD_3 Y10[3] SCLK NET073 S11000X8_LH_YPD_M16
XLH_YPD_2 Y10[2] SCLK NET075 S11000X8_LH_YPD_M16
XLH_YPD_0 Y10[0] SCLK NET070 S11000X8_LH_YPD_M16
XLH_YPD_1 Y10[1] SCLK NET083 S11000X8_LH_YPD_M16
XI154 NET35 Y0N DY[1] S11000X8_SNAND LP2=0.06U WP2=0.18U LP1=0.06U WP1=0.18U LN1=0.06U
+WN1=0.2U LN2=0.06U WN2=0.2U
XI152 NET036 DY[0] Y1N S11000X8_SNAND LP2=0.06U WP2=0.18U LP1=0.06U WP1=0.18U LN1=0.06U
+WN1=0.2U LN2=0.06U WN2=0.2U
XI39 NET41 Y0N Y1N S11000X8_SNAND LP2=0.06U WP2=0.18U LP1=0.06U WP1=0.18U LN1=0.06U WN1=0.2U
+LN2=0.06U WN2=0.2U
XI153 NET53 DY[0] DY[1] S11000X8_SNAND LP2=0.06U WP2=0.18U LP1=0.06U WP1=0.18U LN1=0.06U
+WN1=0.2U LN2=0.06U WN2=0.2U
XI5 DY[0] Y0N S11000X8_SINV LP=0.07U LN=0.07U
XI579 DY[1] Y1N S11000X8_SINV LP=0.07U LN=0.07U
XI200 NET073 NET077 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI199 NET075 NET088 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI123 NET072 NET41 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI124 NET070 NET072 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI202 NET088 NET35 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI190 NET083 NET090 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI201 NET090 NET036 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI215 BISTC BISTT S11000X8_SINV LP=0.07U LN=0.07U
XI203 NET077 NET53 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
**C36 Y1N GND 2F
**C28 DY[0] GND 1.3F
**C27 DY[1] GND 1.3F
**C29 Y0N GND 2F
**C13 NET35 GND 0.5F
**C14 NET088 GND 0.5F
**C15 NET077 GND 0.5F
**C12 NET53 GND 0.5F
**C16 NET090 GND 0.5F
**C17 NET072 GND 0.5F
**C10 NET41 GND 0.5F
**C18 NET070 GND 0.5F
**C19 NET083 GND 0.5F
**C20 NET073 GND 0.5F
**C21 NET075 GND 0.5F
**C11 NET036 GND 0.5F
.ENDS S11000X8_YPRE10_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPREDEC_M16                                                          *
* LAST TIME SAVED: SEP 30 16:22:48 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_YPREDEC_M16 Y10[3] Y10[2] Y10[1] Y10[0] BISTT SCLK Y[1] Y[0] YM[1]
+YM[0]
XYPRE10 Y10[3] Y10[2] Y10[1] Y10[0] BISTT SCLK Y[1] Y[0] YM[1] YM[0] S11000X8_YPRE10_M16
.ENDS S11000X8_YPREDEC_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_XPD8                                                              *
* LAST TIME SAVED: DEC 14 17:25:05 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_LH_XPD8 Q CP D
XI26 NET043 P1 INCPN CP S11000X8_TRANSGATE LP=0.07U WP=3U LN=0.07U WN=1.5U
MN12 GND Q NET39 GND NCH W=0.25U L=0.07U
MN11 NET39 NET042 P1 GND NCH W=0.25U L=0.07U
MP4 NET69 Q VDD VDD PCH W=0.5U L=0.07U
MP5 P1 INCPN NET69 VDD PCH W=0.5U L=0.07U
XI38 NET042 INCPN S11000X8_SINV LP=0.07U WP=0.3U LN=0.07U WN=0.15U
XI24 Q P1 S11000X8_SINV LP=0.07U WP=6U LN=0.07U WN=3U M=2
XI29 INCPN CP S11000X8_SINV LP=0.07U WP=0.5U LN=0.07U WN=0.5U
XI36 NET043 D S11000X8_SINV LP=0.07U WP=3U LN=0.07U WN=1.5U
**C1 INCPN GND 2.759F
**C0 P1 GND 10.654F
**C39 NET042 GND 0.780F
**C3 NET043 GND 3.343F
.ENDS S11000X8_LH_XPD8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XPRE8                                                                *
* LAST TIME SAVED: DEC 14 17:24:55 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_XPRE8 XPRE[7] XPRE[6] XPRE[5] XPRE[4] XPRE[3] XPRE[2] XPRE[1] XPRE[0]
+BIST WLP X[2] X[1] X[0] XM[2] XM[1] XM[0]
MP9 NET51 BISTC X2N VDD PCH W=0.5U L=0.06U
MP0 NET48 BISTC X1N VDD PCH W=0.5U L=0.06U
MP1 VDD X[1] NET39 VDD PCH W=0.5U L=0.06U
MP2 VDD XM[1] NET48 VDD PCH W=0.5U L=0.06U
MP3 NET39 BISTT X1N VDD PCH W=0.5U L=0.06U
MP6 NET36 BISTT X0N VDD PCH W=0.5U L=0.06U
MP7 VDD XM[0] NET27 VDD PCH W=0.5U L=0.06U
MP10 VDD X[0] NET36 VDD PCH W=0.5U L=0.06U
MP11 NET27 BISTC X0N VDD PCH W=0.5U L=0.06U
MP5 VDD X[2] NET60 VDD PCH W=0.5U L=0.06U
MP8 VDD XM[2] NET51 VDD PCH W=0.5U L=0.06U
MP4 NET60 BISTT X2N VDD PCH W=0.5U L=0.06U
MN0 NET84 X[1] GND GND NCH W=0.25U L=0.06U
MN1 NET81 XM[1] GND GND NCH W=0.25U L=0.06U
MN2 X1N BISTC NET84 GND NCH W=0.25U L=0.06U
MN3 X1N BISTT NET81 GND NCH W=0.25U L=0.06U
MN7 NET87 X[2] GND GND NCH W=0.25U L=0.06U
MN8 NET90 XM[2] GND GND NCH W=0.25U L=0.06U
MN4 X2N BISTC NET87 GND NCH W=0.25U L=0.06U
MN6 X0N BISTT NET66 GND NCH W=0.25U L=0.06U
MN9 X0N BISTC NET63 GND NCH W=0.25U L=0.06U
MN10 NET66 XM[0] GND GND NCH W=0.25U L=0.06U
MN11 NET63 X[0] GND GND NCH W=0.25U L=0.06U
MN5 X2N BISTT NET90 GND NCH W=0.25U L=0.06U
XLH_XPD8_2 XPRE[2] WLP NET162 S11000X8_LH_XPD8
XLH_XPD8_3 XPRE[3] WLP NET097 S11000X8_LH_XPD8
XLH_XPD8_7 XPRE[7] WLP NET085 S11000X8_LH_XPD8
XLH_XPD8_5 XPRE[5] WLP NET156 S11000X8_LH_XPD8
XLH_XPD8_1 XPRE[1] WLP NET165 S11000X8_LH_XPD8
XLH_XPD8_6 XPRE[6] WLP NET171 S11000X8_LH_XPD8
XLH_XPD8_0 XPRE[0] WLP NET089 S11000X8_LH_XPD8
XLH_XPD8_4 XPRE[4] WLP NET153 S11000X8_LH_XPD8
XI624 BISTT BISTC S11000X8_SINV LP=0.06U LN=0.06U
XI582 NET165 NET038 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI608 X1 X1N S11000X8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI447 NET089 NET167 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI590 NET156 NET046 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI584 NET097 NET050 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI588 X2 X2N S11000X8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI615 X0 X0N S11000X8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI591 NET171 NET026 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI592 NET085 NET034 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI583 NET162 NET054 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI589 NET153 NET030 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.3U
XI623 BISTC BIST S11000X8_SINV LP=0.06U LN=0.06U
XI600 NET030 X0N X1N X2 S11000X8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI602 NET026 X0N X1 X2 S11000X8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI598 NET054 X0N X1 X2N S11000X8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI603 NET034 X0 X1 X2 S11000X8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI599 NET050 X0 X1 X2N S11000X8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI597 NET038 X0 X1N X2N S11000X8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI407 NET167 X0N X1N X2N S11000X8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
XI601 NET046 X0 X1N X2 S11000X8_SNAND3 LP3=0.06U WP3=0.15U LP2=0.06U WP2=0.15U LP1=0.06U
+WP1=0.15U LN1=0.06U WN1=0.15U LN2=0.06U WN2=0.15U LN3=0.06U WN3=0.15U
**C71 BISTT GND 4.975F
**C72 BISTC GND 5.774F
**C57 NET046 GND 1.321F
**C58 NET030 GND 1.363F
**C67 X1 GND 3.655F
**C68 X1N GND 4.286F
**C66 X2N GND 4.779F
**C46 NET038 GND 1.346F
**C63 NET085 GND 3.233F
**C64 NET156 GND 3.230F
**C65 NET153 GND 3.332F
**C47 NET054 GND 1.329F
**C59 NET165 GND 3.192F
**C50 NET050 GND 1.314F
**C32 X2 GND 3.573F
**C69 X0N GND 6.023F
**C70 X0 GND 5.270F
**C40 NET089 GND 3.244F
**C44 NET167 GND 1.348F
**C60 NET097 GND 3.231F
**C61 NET162 GND 3.239F
**C62 NET171 GND 3.306F
**C55 NET034 GND 1.349F
**C56 NET026 GND 1.307F
.ENDS S11000X8_XPRE8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XPREDEC888                                                           *
* LAST TIME SAVED: DEC  5 14:42:50 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_XPREDEC888 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1]
+XPD0[0] XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0]
+XPD2[7] XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLK
+X[8] X[7] X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4]
+XM[3] XM[2] XM[1] XM[0]
XPRE8_A XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+BIST_BUF SCLK X[2] X[1] X[0] XM[2] XM[1] XM[0] S11000X8_XPRE8
XPRE8_B XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0]
+BIST_BUF SCLK X[5] X[4] X[3] XM[5] XM[4] XM[3] S11000X8_XPRE8
XPRE8_C XPD2[7] XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0]
+BIST_BUF SCLK X[8] X[7] X[6] XM[8] XM[7] XM[6] S11000X8_XPRE8
.ENDS S11000X8_XPREDEC888


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL888_M16                                                          *
* LAST TIME SAVED: DEC  1 14:30:43 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_CTRL888_M16 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7]
+XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2] Y10[1]
+Y10[0] Y32[3] Y32[2] Y32[1] Y32[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1]
+TSEL[0] WEB WEBM WLPTEST X[8] X[7] X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[8]
+XM[7] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0] Y[3] Y[2] Y[1] Y[0] YM[3]
+YM[2] YM[1] YM[0]
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S11000X8_WLPGEN_M16V1
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S11000X8_BISIN_M16
XI180 CTRL_TIEL S11000X8_SRAM_TIEL
XI182 CTRL_TIELB S11000X8_SRAM_TIEL
XYPREDEC32 Y32[3] Y32[2] Y32[1] Y32[0] BIST_BUF NET65 Y[3] Y[2] YM[3] YM[2]
+S11000X8_YPREDEC_M16
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S11000X8_YPREDEC_M16
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[7]
+XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7] XPD2[6]
+XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[8] X[7] X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1]
+XM[0] S11000X8_XPREDEC888
.ENDS S11000X8_CTRL888_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M8V1                                                          *
* LAST TIME SAVED: DEC 14 17:41:43 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_WLPGEN_M8V1 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK TM
+TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 PRE_WLP_RESET D02 SEL[3] SELN[3] SELN[2] S11000X8_DELAY_V3
XI337 D02 PRE_WLP_RESET D01 SEL[2] SELN[2] SELN[1] S11000X8_DELAY_V2
XI326 D01 PRE_WLP_RESET TRWLPBB SEL[1] SELN[1] SELN[0] S11000X8_DELAY_V1
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S11000X8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S11000X8_CLKBUF
XI238 D1 T0 NET259 CLK_K S11000X8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S11000X8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET148 CLK_KB CLK S11000X8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN4 NET151 TRWLPBB GND GND NCH W=0.5U L=0.06U
MN5 PRE_WLP_RESET SEL[0] NET151 GND NCH W=0.5U L=0.06U
MN7 NET165 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET155 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET161 GND NCH W=5U L=0.06U
MN0 NET161 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET165 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET227 NET155 GND NCH W=5U L=0.07U
MP7 NET175 SELN[0] PRE_WLP_RESET VDD PCH W=1.0U L=0.06U
MP10 VDD TRWLPBB NET175 VDD PCH W=1.0U L=0.06U M=1
MP5 VDD TME NET179 VDD PCH W=10U L=0.06U M=2
MP9 NET173 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET186 NET227 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET179 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET173 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET186 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI482 WLP_RESET PRE_WLP_RESET NET217 S11000X8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U
+LN1=0.06U WN1=1.0U LN2=0.06U WN2=1.0U
XI219 NET148 WLP_RESET WLPSTART S11000X8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI328 SELN[0] SEL0N SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S11000X8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI477 NET227 WLPTEST S11000X8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI495 NET209 NET210 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI507 TRWLPBB TRWLPB S11000X8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI494 NET210 NET215 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI386 TRWLPB TRWLP S11000X8_SINV LP=0.12U WP=1.0U LN=0.12U WN=0.4U
XI496 NET218 NET209 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI493 NET215 PRE_WLP_RESET S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI471 SEL[3] SELN[3] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET253 S11000X8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET251 CEB S11000X8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET239 WLPSTART S11000X8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET239 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET243 NET239 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET243 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET239 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI371 NET253 NET251 S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI497 NET217 TRWLP S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI283 CLK_KB CLK S11000X8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
XI296 CLK_K NET259 S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI297 NET259 CLK S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI473 SEL1 SEL1N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI315 TME TMEB S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**C47 SELN[0] GND 2.7F
**C48 SEL[0] GND 2.7F
**C49 SELN[2] GND 2.7F
**C50 SEL[2] GND 2.7F
**C44 SEL[3] GND 2.7F
**C36 TRWLPB GND 5.4F
**C428 D02 GND 1.2F
**C40 NET243 GND 5.6F
**C410 SEL0 GND 2.1F
**C446 TME GND 5.5F
**C426 D01 GND 1.3F
**C420 SEL0N GND 2.9F
**C448 TMEB GND 6.1F
**C0 T2 GND 6.1F
**C4 NET259 GND 0.7F
**C418 SEL1 GND 2.7F
**C34 WLPSTART GND 13.1F
**C35 NET239 GND 8.2F
**C432 NET227 GND 5.2F
**C30 NET253 GND 0.7F
**C43 SELN[3] GND 2.7F
**C29 NET251 GND 0.6F
**C422 SEL1N GND 2.8F
**C32 D1 GND 1.4F
**C1 T1 GND 3.2F
**C5 CLK_K GND 0.8F
**C2 WLP_RESET GND 5.5F
**C430 PRE_WLP_RESET GND 4.2F
**C45 SELN[1] GND 2.7F
**C22 CLK_KB GND 2.2F
**C33 T0 GND 1.0F
**C46 SEL[1] GND 2.7F
**C31 NET148 GND 5.6F
**C51 TRWLPBB GND 5.4F
.ENDS S11000X8_WLPGEN_M8V1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AWTD_M8                                                              *
* LAST TIME SAVED: OCT  4 10:09:37 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_AWTD_M8 AWTI AWT
XINV0 AWTI Z1 S11000X8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI9 Z1 AWT S11000X8_SINV LP=0.07U WP=3U LN=0.07U WN=1.5U
.ENDS S11000X8_AWTD_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISTD_M8                                                             *
* LAST TIME SAVED: OCT  4 10:38:52 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BISTD_M8 BISTC BISTT BIST
XI13 BISTT BISTC S11000X8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI14 BISTC BIST S11000X8_SINV LP=0.07U WP=3.2U LN=0.07U WN=1.6U
.ENDS S11000X8_BISTD_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISIN_M8                                                             *
* LAST TIME SAVED: DEC  1 14:10:29 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BISIN_M8 AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM
XCEBMX CEBX CEB CEBM BISTC BIST_BUF S11000X8_CEBBISMX
XWEBMX WEBX WEB WEBM BISTC BIST_BUF S11000X8_CEBBISMX
XAWTD AWTI AWT S11000X8_AWTD_M8
XBISTD BISTC BIST_BUF BIST S11000X8_BISTD_M8
.ENDS S11000X8_BISIN_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_YPD_M8                                                            *
* LAST TIME SAVED: MAY 25 14:13:06 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_LH_YPD_M8 Q CP D
XI26 D P2 INCPN CP S11000X8_TRANSGATE LP=0.07U WP=2U LN=0.07U WN=2U
MN0 GND Q NET38 GND NCH W=0.2U L=0.07U
MN1 NET38 CP P2 GND NCH W=0.2U L=0.07U
MP4 NET49 Q VDD VDD PCH W=0.5U L=0.07U
MP5 P2 INCPN NET49 VDD PCH W=0.5U L=0.07U
XI23 Q P2 S11000X8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI29 INCPN CP S11000X8_SINV LP=0.07U WP=1.2U LN=0.07U WN=0.6U
**C2 P2 GND 3.9F
**C3 INCPN GND 1.5F
.ENDS S11000X8_LH_YPD_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPRE10_M2                                                            *
* LAST TIME SAVED: SEP 29 14:55:40 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_YPRE10_M2 Y32[1] Y32[0] BISTT SCLK Y[0] YM[0]
MP14 VDD Y[0] Z21 VDD PCH W=0.3U L=0.07U
MP15 Z21 BISTT Y0N VDD PCH W=0.3U L=0.07U
MP7 VDD YM[0] Z22 VDD PCH W=0.3U L=0.07U
MP6 Z22 BISTC Y0N VDD PCH W=0.3U L=0.07U
MN15 Y0N BISTC Z23 GND NCH W=0.15U L=0.07U
MN14 Y0N BISTT Z24 GND NCH W=0.15U L=0.07U
MN6 Z24 YM[0] GND GND NCH W=0.15U L=0.07U
MN13 Z23 Y[0] GND GND NCH W=0.15U L=0.07U
XLH_YPD_0 Y32[0] SCLK NET070 S11000X8_LH_YPD_M8
XLH_YPD_1 Y32[1] SCLK NET083 S11000X8_LH_YPD_M8
XI5 Y0 Y0N S11000X8_SINV LP=0.07U LN=0.07U
XI123 NET072 NET41 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI124 NET070 NET072 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI201 NET083 NET090 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI205 BISTC BISTT S11000X8_SINV LP=0.07U LN=0.07U
XI199 NET41 Y0N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI202 NET090 NET036 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI203 NET036 Y0 S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
**C28 Y0 GND 0.7F
**C29 Y0N GND 1.1F
**C16 NET090 GND 1.1F
**C17 NET072 GND 1.1F
**C10 NET41 GND 1.6F
**C18 NET070 GND 2.9F
**C19 NET083 GND 2.9F
**C11 NET036 GND 1.6F
.ENDS S11000X8_YPRE10_M2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPREDEC_M2                                                           *
* LAST TIME SAVED: OCT 24 09:46:40 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_YPREDEC_M2 Y32[1] Y32[0] BIST_BUF SCLK Y[0] YM[0]
XYPRE10 Y32[1] Y32[0] BIST_BUF SCLK Y[0] YM[0] S11000X8_YPRE10_M2
.ENDS S11000X8_YPREDEC_M2


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPRE10_M8                                                            *
* LAST TIME SAVED: OCT  4 10:00:07 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_YPRE10_M8 Y10[3] Y10[2] Y10[1] Y10[0] BISTT SCLK Y[1] Y[0] YM[1] YM[0]
MN3 Y1N BISTC NET44 GND NCH W=0.15U L=0.07U
MN2 Y1N BISTT NET173 GND NCH W=0.15U L=0.07U
MN15 Y0N BISTC NET174 GND NCH W=0.15U L=0.07U
MN14 Y0N BISTT NET38 GND NCH W=0.15U L=0.07U
MN13 NET174 Y[0] GND GND NCH W=0.15U L=0.07U
MN6 NET38 YM[0] GND GND NCH W=0.15U L=0.07U
MN0 NET173 YM[1] GND GND NCH W=0.15U L=0.07U
MN1 NET44 Y[1] GND GND NCH W=0.15U L=0.07U
MP0 NET47 BISTC Y1N VDD PCH W=0.3U L=0.07U
MP15 NET50 BISTT Y0N VDD PCH W=0.3U L=0.07U
MP14 VDD Y[0] NET50 VDD PCH W=0.3U L=0.07U
MP7 VDD YM[0] NET59 VDD PCH W=0.3U L=0.07U
MP6 NET59 BISTC Y0N VDD PCH W=0.3U L=0.07U
MP1 VDD YM[1] NET47 VDD PCH W=0.3U L=0.07U
MP2 VDD Y[1] NET68 VDD PCH W=0.3U L=0.07U
MP3 NET68 BISTT Y1N VDD PCH W=0.3U L=0.07U
XLH_YPD_3 Y10[3] SCLK NET073 S11000X8_LH_YPD_M8
XLH_YPD_2 Y10[2] SCLK NET075 S11000X8_LH_YPD_M8
XLH_YPD_0 Y10[0] SCLK NET070 S11000X8_LH_YPD_M8
XLH_YPD_1 Y10[1] SCLK NET083 S11000X8_LH_YPD_M8
XI211 NET35 Y0N DY[1] S11000X8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI210 NET036 DY[0] Y1N S11000X8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI212 NET53 DY[0] DY[1] S11000X8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI39 NET41 Y0N Y1N S11000X8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI215 BISTC BISTT S11000X8_SINV LP=0.07U LN=0.07U
XI5 DY[0] Y0N S11000X8_SINV LP=0.07U LN=0.07U
XI579 DY[1] Y1N S11000X8_SINV LP=0.07U LN=0.07U
XI202 NET075 NET088 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI201 NET083 NET090 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI123 NET072 NET41 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI124 NET070 NET072 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI206 NET077 NET53 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI203 NET073 NET077 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI205 NET088 NET35 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI204 NET090 NET036 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
**C36 Y1N GND 2F
**C28 DY[0] GND 1.3F
**C27 DY[1] GND 1.3F
**C29 Y0N GND 2F
**C13 NET35 GND 1.3F
**C14 NET088 GND 1.1F
**C15 NET077 GND 1.1F
**C12 NET53 GND 1.3F
**C16 NET090 GND 1.1F
**C17 NET072 GND 1.1F
**C10 NET41 GND 1.3F
**C18 NET070 GND 2.8F
**C19 NET083 GND 2.8F
**C20 NET073 GND 2.8F
**C21 NET075 GND 2.8F
**C11 NET036 GND 1.3F
.ENDS S11000X8_YPRE10_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPREDEC_M8                                                           *
* LAST TIME SAVED: OCT 24 09:46:40 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_YPREDEC_M8 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF SCLK Y[1] Y[0] YM[1]
+YM[0]
XYPRE10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF SCLK Y[1] Y[0] YM[1] YM[0]
+S11000X8_YPRE10_M8
.ENDS S11000X8_YPREDEC_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL888_M8                                                           *
* LAST TIME SAVED: DEC 14 17:41:45 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_CTRL888_M8 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7]
+XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2] Y10[1]
+Y10[0] Y32[1] Y32[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1] TSEL[0] WEB WEBM
+WLPTEST X[8] X[7] X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5]
+XM[4] XM[3] XM[2] XM[1] XM[0] Y[2] Y[1] Y[0] YM[2] YM[1] YM[0]
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S11000X8_WLPGEN_M8V1
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S11000X8_BISIN_M8
XSRM_TIEL CTRL_TIEL S11000X8_SRAM_TIEL
XSRM_TIEL2 CTRL_TIELB S11000X8_SRAM_TIEL
**C184 SCLKX GND 34.2F
**C187 NET65 GND 15.3F
**C7 WEBX GND 3.022F
XYPREDEC32 Y32[1] Y32[0] BIST_BUF NET65 Y[2] YM[2] S11000X8_YPREDEC_M2
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S11000X8_YPREDEC_M8
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[7]
+XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7] XPD2[6]
+XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[8] X[7] X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1]
+XM[0] S11000X8_XPREDEC888
.ENDS S11000X8_CTRL888_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M4V1                                                          *
* LAST TIME SAVED: DEC 14 16:49:46 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_WLPGEN_M4V1 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK TM
+TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 NET170 D02 SEL[3] SELN[3] SELN[2] S11000X8_DELAY_V3
XI337 D02 NET170 D01 SEL[2] SELN[2] SELN[1] S11000X8_DELAY_V2
XI326 D01 NET170 NET0214 SEL[1] SELN[1] SELN[0] S11000X8_DELAY_V1
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S11000X8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S11000X8_CLKBUF
XI238 D1 T0 NET132 CLK_K S11000X8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S11000X8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET169 CLK_KB CLK S11000X8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN4 NET333 NET0214 GND GND NCH W=0.5U L=0.06U
MN5 NET170 SEL[0] NET333 GND NCH W=0.5U L=0.06U
MN7 NET96 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET097 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET096 GND NCH W=5U L=0.06U
MN0 NET096 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET96 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET0198 NET097 GND NCH W=5U L=0.07U
MP10 VDD NET0214 NET173 VDD PCH W=1.0U L=0.06U M=1
MP5 VDD TME NET0108 VDD PCH W=10U L=0.06U M=2
MP7 NET173 SELN[0] NET170 VDD PCH W=1.0U L=0.06U
MP9 NET80 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET0119 NET0198 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET0108 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET80 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET0119 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI219 NET169 WLP_RESET WLPSTART S11000X8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI482 WLP_RESET NET170 NET218 S11000X8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U LN1=0.06U
+WN1=1.0U LN2=0.06U WN2=1.0U
XI328 SELN[0] SEL0N SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S11000X8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI383 NET0198 WLPTEST S11000X8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI386 TRWLPB TRWLP S11000X8_SINV LP=0.12U WP=1.0U LN=0.12U WN=0.4U
XI496 NET219 NET226 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI494 NET224 NET220 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI471 SEL[3] SELN[3] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET0323 S11000X8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET0321 CEB S11000X8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET0348 WLPSTART S11000X8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET0354 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET0354 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI493 NET220 NET170 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI371 NET0323 NET0321 S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI292 NET0214 TRWLPB S11000X8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI283 CLK_KB CLK S11000X8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
XI296 CLK_K NET132 S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI497 NET218 TRWLP S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI495 NET226 NET224 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI297 NET132 CLK S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI473 SEL1 SEL1N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI315 TME TMEB S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**C36 TRWLPB GND 3.009F
**C44 NET170 GND 5.266F
**C428 D02 GND 1.950F
**C40 NET0354 GND 13.839F
**C43 WLP_RESET GND 4.630F
**C410 SEL0 GND 2.687F
**C446 TME GND 11.753F
**C426 D01 GND 2.319F
**C420 SEL0N GND 2.317F
**C434 NET0214 GND 3.637F
**C448 TMEB GND 11.368F
**C0 T2 GND 9.532F
**C4 NET132 GND 1.008F
**C418 SEL1 GND 2.583F
**C34 WLPSTART GND 28.916F
**C35 NET0348 GND 25.077F
**C432 NET0198 GND 6.135F
**C30 NET0323 GND 1.326F
**C29 NET0321 GND 0.782F
**C422 SEL1N GND 2.592F
**C32 D1 GND 1.821F
**C1 T1 GND 5.899F
**C5 CLK_K GND 1.749F
**C22 CLK_KB GND 6.158F
**C33 T0 GND 3.232F
**C31 NET169 GND 2.156F
.ENDS S11000X8_WLPGEN_M4V1


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: AWTD_M4                                                              *
* LAST TIME SAVED: DEC 14 16:50:10 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_AWTD_M4 AWTI AWT
**C0 Z1 GND 8.034F
XINV0 AWTI Z1 S11000X8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI9 Z1 AWT S11000X8_SINV LP=0.07U WP=3U LN=0.07U WN=1.5U
.ENDS S11000X8_AWTD_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISTD_M4                                                             *
* LAST TIME SAVED: OCT 13 22:07:21 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BISTD_M4 BISTC BIST_BUF BIST
XI13 BIST_BUF BISTC S11000X8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI14 BISTC BIST S11000X8_SINV LP=0.07U WP=3.2U LN=0.07U WN=1.6U
.ENDS S11000X8_BISTD_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BISIN_M4                                                             *
* LAST TIME SAVED: DEC 14 19:54:47 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BISIN_M4 AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM
XCEBMX CEBX CEB CEBM BISTC BIST_BUF S11000X8_CEBBISMX
XWEBMX WEBX WEB WEBM BISTC BIST_BUF S11000X8_CEBBISMX
**C0 BISTC GND 9.597F
XAWTD AWTI AWT S11000X8_AWTD_M4
XBISTD BISTC BIST_BUF BIST S11000X8_BISTD_M4
.ENDS S11000X8_BISIN_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: LH_YPD_M4                                                            *
* LAST TIME SAVED: NOV 10 11:38:58 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_LH_YPD_M4 Q CP D
XI26 D P2 INCPN CP S11000X8_TRANSGATE LP=0.07U WP=2U LN=0.07U WN=2U
MN0 GND Q NET38 GND NCH W=0.2U L=0.07U
MN1 NET38 CP P2 GND NCH W=0.2U L=0.07U
MP4 NET49 Q VDD VDD PCH W=0.5U L=0.07U
MP5 P2 INCPN NET49 VDD PCH W=0.5U L=0.07U
XI23 Q P2 S11000X8_SINV LP=0.07U WP=8U LN=0.07U WN=4U M=2
XI29 INCPN CP S11000X8_SINV LP=0.07U WP=1.2U LN=0.07U WN=0.6U
**C2 P2 GND 13.447F
**C3 INCPN GND 2.178F
.ENDS S11000X8_LH_YPD_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPRE10_M4                                                            *
* LAST TIME SAVED: DEC 14 16:50:11 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_YPRE10_M4 Y10[3] Y10[2] Y10[1] Y10[0] BIST SCLK Y[1] Y[0] YM[1] YM[0]
XLH_YPD_3 Y10[3] SCLK NET073 S11000X8_LH_YPD_M4
XLH_YPD_2 Y10[2] SCLK NET075 S11000X8_LH_YPD_M4
XLH_YPD_0 Y10[0] SCLK NET070 S11000X8_LH_YPD_M4
XLH_YPD_1 Y10[1] SCLK NET083 S11000X8_LH_YPD_M4
MN3 Y1N BISTC NET44 GND NCH W=0.15U L=0.07U
MN2 Y1N BISTT NET173 GND NCH W=0.15U L=0.07U
MN15 Y0N BISTC NET174 GND NCH W=0.15U L=0.07U
MN14 Y0N BISTT NET38 GND NCH W=0.15U L=0.07U
MN13 NET174 Y[0] GND GND NCH W=0.15U L=0.07U
MN6 NET38 YM[0] GND GND NCH W=0.15U L=0.07U
MN0 NET173 YM[1] GND GND NCH W=0.15U L=0.07U
MN1 NET44 Y[1] GND GND NCH W=0.15U L=0.07U
MP0 NET47 BISTC Y1N VDD PCH W=0.3U L=0.07U
MP15 NET50 BISTT Y0N VDD PCH W=0.3U L=0.07U
MP14 VDD Y[0] NET50 VDD PCH W=0.3U L=0.07U
MP7 VDD YM[0] NET59 VDD PCH W=0.3U L=0.07U
MP6 NET59 BISTC Y0N VDD PCH W=0.3U L=0.07U
MP1 VDD YM[1] NET47 VDD PCH W=0.3U L=0.07U
MP2 VDD Y[1] NET68 VDD PCH W=0.3U L=0.07U
MP3 NET68 BISTT Y1N VDD PCH W=0.3U L=0.07U
XI211 NET35 Y0N DY[1] S11000X8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI210 NET036 DY[0] Y1N S11000X8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI212 NET53 DY[0] DY[1] S11000X8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI39 NET41 Y0N Y1N S11000X8_SNAND LP2=0.07U WP2=0.18U LP1=0.07U WP1=0.18U LN1=0.07U
+WN1=0.2U LN2=0.07U WN2=0.2U
XI217 BISTT BISTC S11000X8_SINV LP=0.07U LN=0.07U
XI215 BISTC BIST S11000X8_SINV LP=0.07U LN=0.07U
XI5 DY[0] Y0N S11000X8_SINV LP=0.07U LN=0.07U
XI579 DY[1] Y1N S11000X8_SINV LP=0.07U LN=0.07U
XI202 NET075 NET088 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI201 NET083 NET090 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI123 NET072 NET41 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI124 NET070 NET072 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI206 NET077 NET53 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI203 NET073 NET077 S11000X8_SINV LP=0.07U WP=2U LN=0.07U WN=1U
XI205 NET088 NET35 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
XI204 NET090 NET036 S11000X8_SINV LP=0.07U WP=0.4U LN=0.07U WN=0.2U
**C26 BISTC GND 3.305F
**C30 BISTT GND 2.787F
**C36 Y1N GND 3.008F
**C28 DY[0] GND 1.800F
**C27 DY[1] GND 1.800F
**C29 Y0N GND 3.177F
**C13 NET35 GND 1.134F
**C14 NET088 GND 1.642F
**C15 NET077 GND 1.516F
**C12 NET53 GND 1.460F
**C16 NET090 GND 1.796F
**C17 NET072 GND 1.425F
**C10 NET41 GND 1.330F
**C18 NET070 GND 2.637F
**C19 NET083 GND 2.970F
**C20 NET073 GND 2.854F
**C21 NET075 GND 2.503F
**C11 NET036 GND 1.426F
.ENDS S11000X8_YPRE10_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: YPREDEC_M4                                                           *
* LAST TIME SAVED: OCT 13 22:07:22 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_YPREDEC_M4 Y10[3] Y10[2] Y10[1] Y10[0] BIST SCLK Y[1] Y[0] YM[1] YM[0]
XYPRE10 Y10[3] Y10[2] Y10[1] Y10[0] BIST SCLK Y[1] Y[0] YM[1] YM[0] S11000X8_YPRE10_M4
.ENDS S11000X8_YPREDEC_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL888_M4                                                           *
* LAST TIME SAVED: DEC 14 17:10:45 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_CTRL888_M4 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7]
+XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2] Y10[1]
+Y10[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1] TSEL[0] WEB WEBM WLPTEST X[8]
+X[7] X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4] XM[3]
+XM[2] XM[1] XM[0] Y[1] Y[0] YM[1] YM[0]
**C5 NET241 GND 12.589F
**C6 SCLKX GND 58.558F
**C7 WEBX GND 3.022F
XCTRL_WLPGEN DCLK GW_RB SCLKX NET241 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S11000X8_WLPGEN_M4V1
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S11000X8_BISIN_M4
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET241 Y[1] Y[0] YM[1] YM[0]
+S11000X8_YPREDEC_M4
XI180 CTRL_TIEL S11000X8_SRAM_TIEL
XI182 CTRL_TIELB S11000X8_SRAM_TIEL
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[7]
+XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7] XPD2[6]
+XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[8] X[7] X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[8] XM[7] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1]
+XM[0] S11000X8_XPREDEC888
.ENDS S11000X8_CTRL888_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V6                                                             *
* LAST TIME SAVED: DEC 14 15:09:57 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_DELAY_V6 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET28 TSEL IN S11000X8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI163 OUT_B NET28 S11000X8_SINV_HVT LP=0.16U WP=0.6U LN=0.16U WN=0.3U
**CI153 NET28 GND 0.7F
.ENDS S11000X8_DELAY_V6


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V5                                                             *
* LAST TIME SAVED: DEC 14 15:09:45 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_DELAY_V5 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET44 TSEL IN S11000X8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI165 OUT_B NET44 S11000X8_SINV_HVT LP=0.06U WP=0.6U LN=0.06U WN=0.3U
**CI153 NET44 GND 0.7F
.ENDS S11000X8_DELAY_V5


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: DELAY_V4                                                             *
* LAST TIME SAVED: DEC 15 14:54:17 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_DELAY_V4 OUT_B OUT_A IN SEL SELN TSEL
XI161 NET27 TSEL IN S11000X8_SNAND WP2=0.35U WP1=0.35U WN1=0.35U WN2=0.35U
MN0 OUT_A SEL NET17 GND NCH W=0.5U L=0.06U
MN1 NET17 OUT_B GND GND NCH W=0.5U L=0.06U
MP1 VDD OUT_B NET26 VDD PCH W=1U L=0.06U
MP0 NET26 SELN OUT_A VDD PCH W=1U L=0.06U
XI141 OUT_B NET27 S11000X8_SINV_HVT LP=0.06U WP=0.6U LN=0.06U WN=0.3U
**C151 NET27 GND 0.946F
.ENDS S11000X8_DELAY_V4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M16V3                                                         *
* LAST TIME SAVED: DEC  1 14:40:33 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_WLPGEN_M16V3 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK
+TM TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 NET122 D02 SEL[3] SELN[3] SELN[2] S11000X8_DELAY_V6
XI337 D02 NET122 D01 SEL[2] SELN[2] SELN[1] S11000X8_DELAY_V5
XI326 D01 NET122 NET0214 SEL[1] SELN[1] SELN[0] S11000X8_DELAY_V4
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S11000X8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S11000X8_CLKBUF
**XI324 NET122 NET0214 SEL[0] SELN[0] TRANSGATE LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI324 NET122 NET1227 SEL[0] SELN[0] S11000X8_TRANSGATE LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI238 D1 T0 NET132 CLK_K S11000X8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S11000X8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET169 CLK_KB CLK S11000X8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN7 NET96 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET097 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET096 GND NCH W=5U L=0.06U
MN0 NET096 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET96 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET0198 NET097 GND NCH W=5U L=0.07U
MP5 VDD TME NET0108 VDD PCH W=10U L=0.06U M=2
MP9 NET80 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET0119 NET0198 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET0108 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET80 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET0119 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI219 NET169 WLP_RESET WLPSTART S11000X8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI482 WLP_RESET NET122 NET210 S11000X8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U LN1=0.06U
+WN1=1.0U LN2=0.06U WN2=1.0U
XI328 SELN[0] SEL0N SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S11000X8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI383 NET0198 WLPTEST S11000X8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI386 TRWLPB TRWLP S11000X8_SINV LP=0.2U WP=1.0U LN=0.2U WN=0.4U
XI471 SEL[3] SELN[3] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET0323 S11000X8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET0321 CEB S11000X8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET0348 WLPSTART S11000X8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET0354 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET0354 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI371 NET0323 NET0321 S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI292 NET0214 TRWLPB S11000X8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI283 CLK_KB CLK S11000X8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
**XI493 NET209 NET122 SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI493 NET1227 NET0214 S11000X8_SINV LP=0.06U WP=0.755U LN=0.06U WN=0.2U
XI495 NET213 NET208 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI296 CLK_K NET132 S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI297 NET132 CLK S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**XI494 NET208 NET209 SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI494 NET208 NET122 S11000X8_SINV LP=0.06U WP=0.755U LN=0.06U WN=0.2U
XI473 SEL1 SEL1N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI497 NET210 TRWLP S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI315 TME TMEB S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI496 NET211 NET213 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
**CI414 D03 GND 0.7F
**C36 TRWLPB GND 5.4F
**CI428 D02 GND 1.2F
**C40 NET0354 GND 5.6F
**CI410 SEL0 GND 2.1F
**CI446 TME GND 5.5F
**CI426 D01 GND 1.3F
**CI420 SEL0N GND 2.9F
**CI434 NET0214 GND 1.5F
**CI448 TMEB GND 6.1F
**C0 T2 GND 6.1F
**C4 NET132 GND 0.7F
**CI418 SEL1 GND 2.7F
**C34 WLPSTART GND 13.1F
**C35 NET0348 GND 8.2F
**CI432 NET0198 GND 5.2F
**C30 NET0323 GND 0.7F
**C29 NET0321 GND 0.6F
**CI422 SEL1N GND 2.8F
**C32 D1 GND 1.4F
**C1 T1 GND 3.2F
**C5 CLK_K GND 0.8F
**CI444 SELN[0] GND 3.9F
**C22 CLK_KB GND 2.2F
**CI442 SEL[0] GND 4.1F
**C33 T0 GND 1.0F
**C31 NET169 GND 5.6F
**C2 WLP_RESET GND 5.5F
.ENDS S11000X8_WLPGEN_M16V3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XPRE4                                                                *
* LAST TIME SAVED: DEC 14 15:46:20 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_XPRE4 XPRE[3] XPRE[2] XPRE[1] XPRE[0] BIST WLP X[1] X[0] XM[1] XM[0]
MN11 NET41 X[0] GND GND NCH W=0.25U L=0.06U
MN10 NET38 XM[0] GND GND NCH W=0.25U L=0.06U
MN9 X0N BISTC NET41 GND NCH W=0.25U L=0.06U
MN6 X0N BISTT NET38 GND NCH W=0.25U L=0.06U
MN3 X1N BISTT NET23 GND NCH W=0.25U L=0.06U
MN2 X1N BISTC NET20 GND NCH W=0.25U L=0.06U
MN1 NET23 XM[1] GND GND NCH W=0.25U L=0.06U
MN0 NET20 X[1] GND GND NCH W=0.25U L=0.06U
MP11 NET65 BISTC X0N VDD PCH W=0.5U L=0.06U
MP10 VDD X[0] NET56 VDD PCH W=0.5U L=0.06U
MP7 VDD XM[0] NET65 VDD PCH W=0.5U L=0.06U
MP6 NET56 BISTT X0N VDD PCH W=0.5U L=0.06U
MP3 NET53 BISTT X1N VDD PCH W=0.5U L=0.06U
MP2 VDD XM[1] NET44 VDD PCH W=0.5U L=0.06U
MP1 VDD X[1] NET53 VDD PCH W=0.5U L=0.06U
MP0 NET44 BISTC X1N VDD PCH W=0.5U L=0.06U
XLH_XPD8_2 XPRE[2] WLP NET162 S11000X8_LH_XPD8
XLH_XPD8_3 XPRE[3] WLP NET097 S11000X8_LH_XPD8
XLH_XPD8_1 XPRE[1] WLP NET165 S11000X8_LH_XPD8
XLH_XPD8_0 XPRE[0] WLP NET089 S11000X8_LH_XPD8
XI582 BISTT BISTC S11000X8_SINV LP=0.06U LN=0.06U
XI575 NET165 NET038 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.31U
XI623 BISTC BIST S11000X8_SINV LP=0.06U LN=0.06U
XI615 X0 X0N S11000X8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI608 X1 X1N S11000X8_SINV LP=0.06U WP=0.5U LN=0.06U WN=0.25U
XI447 NET089 NET167 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.31U
XI577 NET097 NET050 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.31U
XI576 NET162 NET054 S11000X8_SINV LP=0.07U WP=0.75U LN=0.07U WN=0.31U
XI574 NET050 X0 X1 S11000X8_SNAND LP2=0.07U WP2=0.15U LP1=0.07U WP1=0.15U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI572 NET038 X0 X1N S11000X8_SNAND LP2=0.07U WP2=0.15U LP1=0.07U WP1=0.15U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI573 NET054 X0N X1 S11000X8_SNAND LP2=0.07U WP2=0.15U LP1=0.07U WP1=0.15U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI407 NET167 X0N X1N S11000X8_SNAND LP2=0.07U WP2=0.15U LP1=0.07U WP1=0.15U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
**C70 X0 GND 1.483F
**C69 X0N GND 3.380F
**C68 X1N GND 2.374F
**C67 X1 GND 1.667F
**C46 NET038 GND 1.453F
**C47 NET054 GND 1.481F
**C59 NET165 GND 3.147F
**C50 NET050 GND 1.384F
**C40 NET089 GND 3.277F
**C44 NET167 GND 1.470F
**C60 NET097 GND 3.216F
**C61 NET162 GND 3.122F
.ENDS S11000X8_XPRE4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: XPREDEC844                                                           *
* LAST TIME SAVED: DEC  6 09:48:41 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_XPREDEC844 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1]
+XPD0[0] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST
+SCLK X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1]
+XM[0]
XPRE4_B XPD1[3] XPD1[2] XPD1[1] XPD1[0] BIST SCLK X[4] X[3] XM[4] XM[3] S11000X8_XPRE4
XPRE4_C XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST SCLK X[6] X[5] XM[6] XM[5] S11000X8_XPRE4
XPRE8_A XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] BIST
+SCLK X[2] X[1] X[0] XM[2] XM[1] XM[0] S11000X8_XPRE8
.ENDS S11000X8_XPREDEC844


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL844_M16                                                          *
* LAST TIME SAVED: DEC  1 14:18:20 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_CTRL844_M16 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2]
+Y10[1] Y10[0] Y32[3] Y32[2] Y32[1] Y32[0] AWT BIST CEB CEBM CLK TM TRWLP
+TSEL[1] TSEL[0] WEB WEBM WLPTEST X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[6]
+XM[5] XM[4] XM[3] XM[2] XM[1] XM[0] Y[3] Y[2] Y[1] Y[0] YM[3] YM[2] YM[1]
+YM[0]
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S11000X8_WLPGEN_M16V3
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S11000X8_BISIN_M16
XI180 CTRL_TIEL S11000X8_SRAM_TIEL
XI182 CTRL_TIELB S11000X8_SRAM_TIEL
XYPREDEC32 Y32[3] Y32[2] Y32[1] Y32[0] BIST_BUF NET65 Y[3] Y[2] YM[3] YM[2]
+S11000X8_YPREDEC_M16
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S11000X8_YPREDEC_M16
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[3]
+XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0]
+S11000X8_XPREDEC844
.ENDS S11000X8_CTRL844_M16


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M8V3                                                          *
* LAST TIME SAVED: DEC 14 19:38:34 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_WLPGEN_M8V3 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK TM
+TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 PRE_WLP_RESET D02 SEL[3] SELN[3] SELN[2] S11000X8_DELAY_V6
XI337 D02 PRE_WLP_RESET D01 SEL[2] SELN[2] SELN[1] S11000X8_DELAY_V5
XI326 D01 PRE_WLP_RESET TRWLPBB SEL[1] SELN[1] SELN[0] S11000X8_DELAY_V4
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S11000X8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S11000X8_CLKBUF
XI238 D1 T0 NET259 CLK_K S11000X8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S11000X8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET148 CLK_KB CLK S11000X8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN4 NET151 TRWLPBB GND GND NCH W=0.5U L=0.06U
MN5 PRE_WLP_RESET SEL[0] NET151 GND NCH W=0.5U L=0.06U
MN7 NET165 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET155 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET161 GND NCH W=5U L=0.06U
MN0 NET161 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET165 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET227 NET155 GND NCH W=5U L=0.07U
MP7 NET175 SELN[0] PRE_WLP_RESET VDD PCH W=1.0U L=0.06U
MP10 VDD TRWLPBB NET175 VDD PCH W=1.0U L=0.06U M=1
MP5 VDD TME NET179 VDD PCH W=10U L=0.06U M=2
MP9 NET173 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET186 NET227 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET179 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET173 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET186 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI482 WLP_RESET PRE_WLP_RESET NET217 S11000X8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U
+LN1=0.06U WN1=1.0U LN2=0.06U WN2=1.0U
XI219 NET148 WLP_RESET WLPSTART S11000X8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI328 SELN[0] SEL0N SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S11000X8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI477 NET227 WLPTEST S11000X8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI495 NET209 NET210 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI507 TRWLPBB TRWLPB S11000X8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI494 NET210 NET215 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI386 TRWLPB TRWLP S11000X8_SINV LP=0.12U WP=1.0U LN=0.12U WN=0.4U
XI496 NET218 NET209 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI493 NET215 PRE_WLP_RESET S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI471 SEL[3] SELN[3] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET253 S11000X8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET251 CEB S11000X8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET239 WLPSTART S11000X8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET239 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET243 NET239 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET243 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET239 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI371 NET253 NET251 S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI497 NET217 TRWLP S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI283 CLK_KB CLK S11000X8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
XI296 CLK_K NET259 S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI297 NET259 CLK S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI473 SEL1 SEL1N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI315 TME TMEB S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**C47 SELN[0] GND 2.7F
**C48 SEL[0] GND 2.7F
**C49 SELN[2] GND 2.7F
**C50 SEL[2] GND 2.7F
**C44 SEL[3] GND 2.7F
**C36 TRWLPB GND 5.4F
**CI428 D02 GND 1.2F
**C40 NET243 GND 5.6F
**CI410 SEL0 GND 2.1F
**CI446 TME GND 5.5F
**CI426 D01 GND 1.3F
**CI420 SEL0N GND 2.9F
**CI448 TMEB GND 6.1F
**C0 T2 GND 6.1F
**C4 NET259 GND 0.7F
**CI418 SEL1 GND 2.7F
**C34 WLPSTART GND 13.1F
**C35 NET239 GND 8.2F
**CI432 NET227 GND 5.2F
**C30 NET253 GND 0.7F
**C43 SELN[3] GND 2.7F
**C15 NET251 GND 0.7F
**CI422 SEL1N GND 2.8F
**C32 D1 GND 1.4F
**C1 T1 GND 3.2F
**C5 CLK_K GND 0.8F
**C2 WLP_RESET GND 5.5F
**CI430 PRE_WLP_RESET GND 4.2F
**C45 SELN[1] GND 2.7F
**C22 CLK_KB GND 2.2F
**C33 T0 GND 1.0F
**C46 SEL[1] GND 2.7F
**C31 NET148 GND 5.6F
**C51 TRWLPBB GND 5.4F
.ENDS S11000X8_WLPGEN_M8V3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL844_M8                                                           *
* LAST TIME SAVED: DEC 14 19:38:13 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_CTRL844_M8 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2]
+Y10[1] Y10[0] Y32[1] Y32[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1] TSEL[0] WEB
+WEBM WLPTEST X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2]
+XM[1] XM[0] Y[2] Y[1] Y[0] YM[2] YM[1] YM[0]
**C16 BIST_BUF GND 29.489F
**C5 NET65 GND 12.844F
**C6 SCLKX GND 42.727F
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S11000X8_WLPGEN_M8V3
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S11000X8_BISIN_M8
XI180 CTRL_TIEL S11000X8_SRAM_TIEL
XI182 CTRL_TIELB S11000X8_SRAM_TIEL
XYPREDEC32 Y32[1] Y32[0] BIST_BUF NET65 Y[2] YM[2] S11000X8_YPREDEC_M2
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S11000X8_YPREDEC_M8
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[3]
+XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0]
+S11000X8_XPREDEC844
.ENDS S11000X8_CTRL844_M8


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: WLPGEN_M4V3                                                          *
* LAST TIME SAVED: DEC 14 16:35:44 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_WLPGEN_M4V3 DCLK GW_RB SCLK_X SCLK_Y WLPX WLPY WLPYB0 WLPYB1 CEB CLK TM
+TRWLP TSEL[1] TSEL[0] WEB WLPTEST
XI339 D03 NET170 D02 SEL[3] SELN[3] SELN[2] S11000X8_DELAY_V6
XI337 D02 NET170 D01 SEL[2] SELN[2] SELN[1] S11000X8_DELAY_V5
XI326 D01 NET170 NET0214 SEL[1] SELN[1] SELN[0] S11000X8_DELAY_V4
XPREBUF SCLK_X SCLK_Y CEB CLK WLPX S11000X8_PREBUF
XCLKBUF DCLK GW_RB CEB CLK WEB S11000X8_CLKBUF
XI238 D1 T0 NET132 CLK_K S11000X8_TRANSGATE LP=0.06U WP=1U LN=0.06U WN=0.5U
XI228 T1 T2 CLK CLK_KB S11000X8_TRANSGATE LP=0.06U WP=6U LN=0.06U WN=3U
XI100 T2 NET169 CLK_KB CLK S11000X8_TRANSGATE LP=0.06U WP=1.6U LN=0.06U WN=0.8U
MN4 NET333 NET0214 GND GND NCH W=0.5U L=0.06U
MN5 NET170 SEL[0] NET333 GND NCH W=0.5U L=0.06U
MN7 NET96 CLK_K T0 GND NCH W=0.3U L=0.06U
MN3 NET097 TME GND GND NCH W=10U L=0.07U
MN1 WLPSTART T2 NET096 GND NCH W=5U L=0.06U
MN0 NET096 TMEB GND GND NCH W=8U L=0.06U
MN8 GND T1 NET96 GND NCH W=0.3U L=0.06U
MN2 WLPSTART NET0198 NET097 GND NCH W=5U L=0.07U
MP10 VDD NET0214 NET173 VDD PCH W=1.0U L=0.06U M=1
MP5 VDD TME NET0108 VDD PCH W=10U L=0.06U M=2
MP7 NET173 SELN[0] NET170 VDD PCH W=1.0U L=0.06U
MP9 NET80 T1 VDD VDD PCH W=0.6U L=0.06U
MP2 NET0119 NET0198 WLPSTART VDD PCH W=10U L=0.07U
MP1 NET0108 T2 WLPSTART VDD PCH W=6U L=0.06U M=2
MP8 T0 CLK_KB NET80 VDD PCH W=0.6U L=0.06U
MP3 VDD TMEB NET0119 VDD PCH W=10U L=0.07U M=2
XI468 SELN[3] SEL0 SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI219 NET169 WLP_RESET WLPSTART S11000X8_SNAND LP2=0.06U WP2=1.6U LP1=0.06U WP1=1.6U
+LN1=0.06U WN1=0.8U LN2=0.06U WN2=0.8U
XI482 WLP_RESET NET170 NET218 S11000X8_SNAND LP2=0.06U WP2=1.0U LP1=0.06U WP1=1.0U LN1=0.06U
+WN1=1.0U LN2=0.06U WN2=1.0U
XI328 SELN[0] SEL0N SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI467 SELN[2] SEL0N SEL1 S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI466 SELN[1] SEL0 SEL1N S11000X8_SNAND LP2=0.07U WP2=0.2U LP1=0.07U WP1=0.2U LN1=0.07U
+WN1=0.15U LN2=0.07U WN2=0.15U
XI237 T1 WLP_RESET T0 S11000X8_SNAND LP2=0.06U WP2=3U LP1=0.06U WP1=3U LN1=0.06U WN1=2U
+LN2=0.06U WN2=2U
XI383 NET0198 WLPTEST S11000X8_SINV LP=0.07U WP=4U LN=0.07U WN=2U
XI386 TRWLPB TRWLP S11000X8_SINV LP=0.12U WP=1.0U LN=0.12U WN=0.4U
XI496 NET219 NET226 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI494 NET224 NET220 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI471 SEL[3] SELN[3] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI199 D1 NET0323 S11000X8_SINV LP=0.06U WP=1.2U LN=0.06U WN=0.6U
XI266 NET0321 CEB S11000X8_SINV LP=0.10U WP=0.30U LN=0.10U WN=0.15U
XI308 SEL0N TSEL[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI166 NET0348 WLPSTART S11000X8_SINV LP=0.06U WP=6U LN=0.06U WN=6U M=2
XI156 WLPYB1 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI171 NET0354 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U
XI157 WLPY NET0354 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI168 WLPYB0 NET0348 S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=4U M=2
XI164 WLPX WLPSTART S11000X8_SINV LP=0.06U WP=10U LN=0.06U WN=10U M=2
XI493 NET220 NET170 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI371 NET0323 NET0321 S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI292 NET0214 TRWLPB S11000X8_SINV LP=0.06U WP=1.0U LN=0.06U WN=0.5U
XI283 CLK_KB CLK S11000X8_SINV LP=0.06U WP=2U LN=0.06U WN=1U
XI296 CLK_K NET132 S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI497 NET218 TRWLP S11000X8_SINV LP=0.06U WP=0.4U LN=0.06U WN=0.2U
XI495 NET226 NET224 S11000X8_SINV LP=0.24U WP=0.4U LN=0.24U WN=0.2U
XI297 NET132 CLK S11000X8_SINV LP=0.06U WP=0.6U LN=0.06U WN=0.3U
XI317 TMEB TM S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
XI473 SEL1 SEL1N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI452 SEL0 SEL0N S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI470 SEL[2] SELN[2] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI472 SEL1N TSEL[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI332 SEL[0] SELN[0] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI469 SEL[1] SELN[1] S11000X8_SINV LP=0.07U WP=0.28U LN=0.07U WN=0.15U
XI315 TME TMEB S11000X8_SINV LP=0.07U WP=1U LN=0.07U WN=0.5U
**C36 TRWLPB GND 3.301F
**C428 D02 GND 1.848F
**C40 NET0354 GND 13.287F
**C43 WLP_RESET GND 4.827F
**C410 SEL0 GND 2.559F
**C446 TME GND 11.593F
**C426 D01 GND 2.144F
**C420 SEL0N GND 2.663F
**C434 NET0214 GND 3.842F
**C448 TMEB GND 11.386F
**C0 T2 GND 10.101F
**C4 NET132 GND 0.992F
**C418 SEL1 GND 2.410F
**C34 WLPSTART GND 29.449F
**C35 NET0348 GND 25.222F
**CI432 NET0198 GND 5.2F
**C30 NET0323 GND 1.156F
**C15 NET0321 GND 0.780F
**C422 SEL1N GND 2.768F
**C32 D1 GND 1.699F
**C1 T1 GND 5.839F
**C5 CLK_K GND 1.716F
**C22 CLK_KB GND 6.404F
**C33 T0 GND 3.299F
**C31 NET169 GND 2.481F
.ENDS S11000X8_WLPGEN_M4V3


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CTRL844_M4                                                           *
* LAST TIME SAVED: DEC 14 15:38:03 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_CTRL844_M4 AWTI BIST_BUF CTRL_TIEL CTRL_TIELB DCLK GW_RB WLPX WLPY
+WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0]
+XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2]
+Y10[1] Y10[0] AWT BIST CEB CEBM CLK TM TRWLP TSEL[1] TSEL[0] WEB WEBM WLPTEST
+X[6] X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0]
+Y[1] Y[0] YM[1] YM[0]
**C7 WEBX GND 2.856F
**C16 BIST_BUF GND 29.489F
**C6 SCLKX GND 42.727F
**C5 NET65 GND 12.844F
XCTRL_WLPGEN DCLK GW_RB SCLKX NET65 WLPX WLPY WLPYB0 WLPYB1 CEBX CLK TM TRWLP
+TSEL[1] TSEL[0] WEBX WLPTEST S11000X8_WLPGEN_M4V3
XBIST AWTI BIST_BUF CEBX WEBX AWT BIST CEB CEBM WEB WEBM S11000X8_BISIN_M4
XYPREDEC10 Y10[3] Y10[2] Y10[1] Y10[0] BIST_BUF NET65 Y[1] Y[0] YM[1] YM[0]
+S11000X8_YPREDEC_M4
XI180 CTRL_TIEL S11000X8_SRAM_TIEL
XI182 CTRL_TIELB S11000X8_SRAM_TIEL
XPREDEC XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[3]
+XPD1[2] XPD1[1] XPD1[0] XPD2[3] XPD2[2] XPD2[1] XPD2[0] BIST_BUF SCLKX X[6]
+X[5] X[4] X[3] X[2] X[1] X[0] XM[6] XM[5] XM[4] XM[3] XM[2] XM[1] XM[0]
+S11000X8_XPREDEC844
.ENDS S11000X8_CTRL844_M4


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: MDEC_TRK                                                             *
* LAST TIME SAVED: DEC 14 16:50:12 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_MDEC_TRK WLOUT WLPY WLPYB
XI280 WLOUT NET21 S11000X8_SINV_HVTP LN=0.06U WN=5U    LP=0.07U WP=10U    M=2
XI290 NET33 NET15 S11000X8_SINV LP=0.06U WP=0.8U  LN=0.06U WN=0.8U 
MN2 NET15 NET25 GND GND NCH W=0.5U L=0.06U
MN0 NET21 NET33 WLPY GND NCH W=2.0U   L=0.06U
MN1 NET20 NET20 GND GND NCH W=0.5U L=0.06U
MP0 VDD NET33 NET21 VDD PCH W=2.0U   L=0.06U
MP1 NET21 WLPYB VDD VDD PCH W=2.0U      L=0.06U
MP2 VDD NET20 NET25 VDD PCH W=1U L=0.06U
**C3 NET21 GND 9.553F
**C4 NET33 GND 3.064F
.ENDS S11000X8_MDEC_TRK


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: BCELL                                                                *
* LAST TIME SAVED: OCT 19 14:40:20 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_BCELL BL BLB WL
MN1 BL_IN BLB_IN GND GND NCHPD_HVTSR W=0.14U  L=0.065U  AD=0.02P AS=0.011P PD=0.6U
+PS=0.3U
MN5 GND BL_IN BLB_IN GND NCHPD_HVTSR W=0.14U  L=0.065U  AD=0.02P AS=0.011P PD=0.6U
+PS=0.3U
MN3 BL WL BL_IN GND NCHPG_HVTSR W=0.09U  L=0.075U AD=0.02P AS=0.008P PD=0.6U PS=0.275U
MN0 BLB_IN WL BLB GND NCHPG_HVTSR W=0.09U  L=0.075U AD=0.02P AS=0.008P PD=0.6U
+PS=0.275U
MP2 VDD BL_IN BLB_IN VDD PCHPU_HVTSR W=0.08U  L=0.065U  AD=0.009P AS=0.008P PD=0.34U
+PS=0.265U
MP0 BL_IN BLB_IN VDD VDD PCHPU_HVTSR W=0.08U  L=0.065U  AD=0.009P AS=0.008P PD=0.34U
+PS=0.265U
**C1 BL_IN GND 0.15F
**C0 BLB_IN GND 0.15F
.ENDS S11000X8_BCELL


*******************************************************************************
* SUB-CIRCUIT NETLIST:                                                        *
*                                                                             *
* BLOCK: CELLX4                                                               *
* LAST TIME SAVED: MAY 17 15:57:24 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_CELLX4 BL[0] BL[1] BLB[0] BLB[1] WL[0] WL[1]
XI7 BLB[1] BL[1] WL[1] S11000X8_BCELL
XBCELL1 BLB[1] BL[1] WL[0] S11000X8_BCELL
XI6 BLB[0] BL[0] WL[1] S11000X8_BCELL
XBCELL0 BLB[0] BL[0] WL[0] S11000X8_BCELL
.ENDS S11000X8_CELLX4


*******************************************************************************
* MAIN CIRCUIT NETLIST:                                                       *
*                                                                             *
* BLOCK: LEAFCELL                                                             *
* LAST TIME SAVED: DEC 15 15:43:07 2005                                       *
*******************************************************************************
.SUBCKT S11000X8_LEAFCELL
XI25 NET183[0] NET183[1] NET184 NET185 NET182[0] NET182[1] S11000X8_TRKDUMX2
XI24 NET187[0] NET187[1] NET189 NET190 NET188 NET186[0] NET186[1] S11000X8_TRKNORX2
XI23 NET192[0] NET192[1] NET101 NET195 NET193 NET191[0] NET191[1] S11000X8_TRKMINX2
XI3 NET11 NET412 NET486 NET8 NET7 S11000X8_TRKMIN
XI4 NET6 NET4 NET459 NET13 NET22 NET23 S11000X8_TRKNOR
XI2 NET17 NET15 NET492 NET442 NET12 S11000X8_TRKDUM
XI21 NET473 S11000X8_SRAM_TIEH
XI17 NET0306[0] NET0306[1] NET0306[2] NET0306[3] NET268 NET315 NET260
+NET0305[0] NET0305[1] NET0305[2] NET0305[3] NET312 NET281 S11000X8_XDRVX2
XI8 NET155 NET147[0] NET147[1] NET147[2] NET147[3] NET147[4] NET147[5]
+NET147[6] NET147[7] NET147[8] NET147[9] NET147[10] NET147[11] NET147[12]
+NET147[13] NET147[14] NET147[15] NET146[0] NET146[1] NET146[2] NET146[3]
+NET146[4] NET146[5] NET146[6] NET146[7] NET146[8] NET146[9] NET146[10]
+NET146[11] NET146[12] NET146[13] NET146[14] NET146[15] NET254 NET330 NET154
+NET252 NET153 NET152 NET253 NET151 NET149 NET148[0] NET148[1] NET148[2]
+NET148[3] NET145[0] NET145[1] NET145[2] NET145[3] S11000X8_IO_M16
XI7 NET166 NET156[0] NET156[1] NET156[2] NET156[3] NET156[4] NET156[5]
+NET156[6] NET156[7] NET157[0] NET157[1] NET157[2] NET157[3] NET157[4]
+NET157[5] NET157[6] NET157[7] NET269 NET221 NET165 NET267 NET164 NET163 NET266
+NET162 NET160 NET159[0] NET159[1] NET159[2] NET159[3] NET158[0] NET158[1]
+S11000X8_IO_M8
XI6 NET174 NET175[0] NET175[1] NET175[2] NET175[3] NET176[0] NET176[1]
+NET176[2] NET176[3] NET280 NET194 NET173 NET282 NET172 NET171 NET45 NET170
+NET168 NET167[0] NET167[1] NET167[2] NET167[3] S11000X8_IO_M4
XI14 NET300 NET334 NET381 NET229 NET216 NET213 NET20 NET19 NET18 NET203
+NET207[0] NET207[1] NET207[2] NET207[3] NET207[4] NET207[5] NET207[6]
+NET207[7] NET325[0] NET325[1] NET325[2] NET325[3] NET325[4] NET325[5]
+NET325[6] NET325[7] NET326[0] NET326[1] NET326[2] NET326[3] NET326[4]
+NET326[5] NET326[6] NET326[7] NET208[0] NET208[1] NET208[2] NET208[3]
+NET214[0] NET214[1] NET214[2] NET214[3] NET296 NET295 NET223 NET299 NET201
+NET224 NET217 NET211[0] NET211[1] NET220 NET294 NET112 NET324[0] NET324[1]
+NET324[2] NET324[3] NET324[4] NET324[5] NET324[6] NET324[7] NET324[8]
+NET293[0] NET293[1] NET293[2] NET293[3] NET293[4] NET293[5] NET293[6]
+NET293[7] NET293[8] NET219[0] NET219[1] NET219[2] NET219[3] NET297[0]
+NET297[1] NET297[2] NET297[3] S11000X8_CTRL888_M16
XI13 NET331 NET144 NET405 NET415 NET72 NET71 NET69 NET68 NET67 NET66 NET65[0]
+NET65[1] NET65[2] NET65[3] NET65[4] NET65[5] NET65[6] NET65[7] NET349[0]
+NET349[1] NET349[2] NET349[3] NET349[4] NET349[5] NET349[6] NET349[7]
+NET350[0] NET350[1] NET350[2] NET350[3] NET350[4] NET350[5] NET350[6]
+NET350[7] NET62[0] NET62[1] NET62[2] NET62[3] NET51[0] NET51[1] NET64 NET70
+NET61 NET328 NET60 NET58 NET57 NET56[0] NET56[1] NET55 NET327 NET233 NET348[0]
+NET348[1] NET348[2] NET348[3] NET348[4] NET348[5] NET348[6] NET348[7]
+NET348[8] NET332[0] NET332[1] NET332[2] NET332[3] NET332[4] NET332[5]
+NET332[6] NET332[7] NET332[8] NET49[0] NET49[1] NET49[2] NET333[0] NET333[1]
+NET333[2] S11000X8_CTRL888_M8
XI12 NET364 NET234 NET431 NET401 NET120 NET119 NET117 NET116 NET115 NET114
+NET113[0] NET113[1] NET113[2] NET113[3] NET113[4] NET113[5] NET113[6]
+NET113[7] NET375[0] NET375[1] NET375[2] NET375[3] NET375[4] NET375[5]
+NET375[6] NET375[7] NET374[0] NET374[1] NET374[2] NET374[3] NET374[4]
+NET374[5] NET374[6] NET374[7] NET110[0] NET110[1] NET110[2] NET110[3] NET362
+NET363 NET109 NET359 NET108 NET106 NET105 NET104[0] NET104[1] NET103 NET357
+NET205 NET373[0] NET373[1] NET373[2] NET373[3] NET373[4] NET373[5] NET373[6]
+NET373[7] NET373[8] NET360[0] NET360[1] NET360[2] NET360[3] NET360[4]
+NET360[5] NET360[6] NET360[7] NET360[8] NET99[0] NET99[1] NET361[0] NET361[1]
+S11000X8_CTRL888_M4
XI11 NET395 NET414 NET455 NET413 NET47 NET46 NET44 NET43 NET42 NET41 NET40[0]
+NET40[1] NET40[2] NET40[3] NET40[4] NET40[5] NET40[6] NET40[7] NET39[0]
+NET39[1] NET39[2] NET39[3] NET38[0] NET38[1] NET38[2] NET38[3] NET37[0]
+NET37[1] NET37[2] NET37[3] NET26[0] NET26[1] NET26[2] NET26[3] NET394 NET393
+NET206 NET389 NET222 NET204 NET32 NET31[0] NET31[1] NET30 NET390 NET231
+NET27[0] NET27[1] NET27[2] NET27[3] NET27[4] NET27[5] NET27[6] NET391[0]
+NET391[1] NET391[2] NET391[3] NET391[4] NET391[5] NET391[6] NET25[0] NET25[1]
+NET25[2] NET25[3] NET392[0] NET392[1] NET392[2] NET392[3] S11000X8_CTRL844_M16
XI10 NET428 NET444 NET479 NET445 NET97 NET96 NET94 NET93 NET92 NET91 NET90[0]
+NET90[1] NET90[2] NET90[3] NET90[4] NET90[5] NET90[6] NET90[7] NET89[0]
+NET89[1] NET89[2] NET89[3] NET88[0] NET88[1] NET88[2] NET88[3] NET87[0]
+NET87[1] NET87[2] NET87[3] NET76[0] NET76[1] NET421 NET420 NET86 NET426 NET85
+NET83 NET82 NET81[0] NET81[1] NET80 NET424 NET235 NET77[0] NET77[1] NET77[2]
+NET77[3] NET77[4] NET77[5] NET77[6] NET423[0] NET423[1] NET423[2] NET423[3]
+NET423[4] NET423[5] NET423[6] NET74[0] NET74[1] NET74[2] NET422[0] NET422[1]
+NET422[2] S11000X8_CTRL844_M8
XI9 NET460 NET236 NET505 NET475 NET143 NET142 NET140 NET139 NET138 NET137
+NET136[0] NET136[1] NET136[2] NET136[3] NET136[4] NET136[5] NET136[6]
+NET136[7] NET135[0] NET135[1] NET135[2] NET135[3] NET134[0] NET134[1]
+NET134[2] NET134[3] NET133[0] NET133[1] NET133[2] NET133[3] NET458 NET457
+NET132 NET453 NET131 NET129 NET128 NET127[0] NET127[1] NET126 NET48 NET84
+NET123[0] NET123[1] NET123[2] NET123[3] NET123[4] NET123[5] NET123[6] NET52[0]
+NET52[1] NET52[2] NET52[3] NET52[4] NET52[5] NET52[6] NET122[0] NET122[1]
+NET456[0] NET456[1] S11000X8_CTRL844_M4
XI16 NET227 NET226 NET225 S11000X8_MDEC_TRK
XI1 NET3[0] NET3[1] NET2[0] NET2[1] NET1[0] NET1[1] S11000X8_CELLX4
D7 GND NET322 NDIO W=1.2U L=1.8U
.ENDS S11000X8_LEAFCELL


**** End of leaf cells

.SUBCKT S11000X8_DECODER TRKBL TIEH WL[511] WL[510] WL[509] WL[508] WL[507] 
+ WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] 
+ WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] 
+ WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] 
+ WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] 
+ WL[470] WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] 
+ WL[461] WL[460] WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] 
+ WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] 
+ WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436] WL[435] 
+ WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426] 
+ WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] 
+ WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] 
+ WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] 
+ WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] 
+ WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] 
+ WL[380] WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] 
+ WL[371] WL[370] WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] 
+ WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] 
+ WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346] WL[345] 
+ WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336] 
+ WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] 
+ WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] 
+ WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] 
+ WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] 
+ WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] 
+ WL[290] WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] 
+ WL[281] WL[280] WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] 
+ WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] 
+ WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256] WL[255] 
+ WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] 
+ WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] 
+ WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] 
+ WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] 
+ WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] 
+ WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] 
+ WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] 
+ WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] 
+ WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] 
+ WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] 
+ WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] 
+ WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] 
+ WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] 
+ WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] 
+ WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] 
+ WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] 
+ WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] 
+ WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] 
+ WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] 
+ WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] 
+ WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] 
+ WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] 
+ WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] 
+ WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] 
+ WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] 
+ WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] 
+ WL[2] WL[1] WL[0] TRKWL WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] 
+ XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] 
+ XPD1[2] XPD1[1] XPD1[0] XPD2[7] XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] 
+ XPD2[1] XPD2[0]
XTIEH TIEH S11000X8_SRAM_TIEH
XDECTRK TRKWL WLPY WLPYB0 S11000X8_MDEC_TRK
MP1 VDD TRKWL TRKBL VDD PCH W=2.1U L=0.07U
XDEC0 WL[1] WL[0] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[0]
+  S11000X8_XDRV
XDEC1 WL[2] WL[3] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[0]
+  S11000X8_XDRV
XDEC2 WL[5] WL[4] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[0]
+  S11000X8_XDRV
XDEC3 WL[6] WL[7] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[0]
+  S11000X8_XDRV
XDEC4 WL[9] WL[8] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[0]
+  S11000X8_XDRV
XDEC5 WL[10] WL[11] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[0]
+  S11000X8_XDRV
XDEC6 WL[13] WL[12] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[0]
+  S11000X8_XDRV
XDEC7 WL[14] WL[15] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[0]
+  S11000X8_XDRV
XDEC8 WL[17] WL[16] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[0]
+  S11000X8_XDRV
XDEC9 WL[18] WL[19] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[0]
+  S11000X8_XDRV
XDEC10 WL[21] WL[20] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[0]
+  S11000X8_XDRV
XDEC11 WL[22] WL[23] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[0]
+  S11000X8_XDRV
XDEC12 WL[25] WL[24] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[0]
+  S11000X8_XDRV
XDEC13 WL[26] WL[27] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[0]
+  S11000X8_XDRV
XDEC14 WL[29] WL[28] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[0]
+  S11000X8_XDRV
XDEC15 WL[30] WL[31] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[0]
+  S11000X8_XDRV
XDEC16 WL[33] WL[32] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[4] XPD2[0]
+  S11000X8_XDRV
XDEC17 WL[34] WL[35] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[4] XPD2[0]
+  S11000X8_XDRV
XDEC18 WL[37] WL[36] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[4] XPD2[0]
+  S11000X8_XDRV
XDEC19 WL[38] WL[39] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[4] XPD2[0]
+  S11000X8_XDRV
XDEC20 WL[41] WL[40] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[5] XPD2[0]
+  S11000X8_XDRV
XDEC21 WL[42] WL[43] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[5] XPD2[0]
+  S11000X8_XDRV
XDEC22 WL[45] WL[44] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[5] XPD2[0]
+  S11000X8_XDRV
XDEC23 WL[46] WL[47] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[5] XPD2[0]
+  S11000X8_XDRV
XDEC24 WL[49] WL[48] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[6] XPD2[0]
+  S11000X8_XDRV
XDEC25 WL[50] WL[51] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[6] XPD2[0]
+  S11000X8_XDRV
XDEC26 WL[53] WL[52] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[6] XPD2[0]
+  S11000X8_XDRV
XDEC27 WL[54] WL[55] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[6] XPD2[0]
+  S11000X8_XDRV
XDEC28 WL[57] WL[56] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[7] XPD2[0]
+  S11000X8_XDRV
XDEC29 WL[58] WL[59] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[7] XPD2[0]
+  S11000X8_XDRV
XDEC30 WL[61] WL[60] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[7] XPD2[0]
+  S11000X8_XDRV
XDEC31 WL[62] WL[63] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[7] XPD2[0]
+  S11000X8_XDRV
XDEC32 WL[65] WL[64] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[1]
+  S11000X8_XDRV
XDEC33 WL[66] WL[67] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[1]
+  S11000X8_XDRV
XDEC34 WL[69] WL[68] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[1]
+  S11000X8_XDRV
XDEC35 WL[70] WL[71] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[1]
+  S11000X8_XDRV
XDEC36 WL[73] WL[72] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[1]
+  S11000X8_XDRV
XDEC37 WL[74] WL[75] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[1]
+  S11000X8_XDRV
XDEC38 WL[77] WL[76] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[1]
+  S11000X8_XDRV
XDEC39 WL[78] WL[79] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[1]
+  S11000X8_XDRV
XDEC40 WL[81] WL[80] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[1]
+  S11000X8_XDRV
XDEC41 WL[82] WL[83] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[1]
+  S11000X8_XDRV
XDEC42 WL[85] WL[84] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[1]
+  S11000X8_XDRV
XDEC43 WL[86] WL[87] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[1]
+  S11000X8_XDRV
XDEC44 WL[89] WL[88] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[1]
+  S11000X8_XDRV
XDEC45 WL[90] WL[91] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[1]
+  S11000X8_XDRV
XDEC46 WL[93] WL[92] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[1]
+  S11000X8_XDRV
XDEC47 WL[94] WL[95] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[1]
+  S11000X8_XDRV
XDEC48 WL[97] WL[96] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[4] XPD2[1]
+  S11000X8_XDRV
XDEC49 WL[98] WL[99] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[4] XPD2[1]
+  S11000X8_XDRV
XDEC50 WL[101] WL[100] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[4] XPD2[1]
+  S11000X8_XDRV
XDEC51 WL[102] WL[103] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[4] XPD2[1]
+  S11000X8_XDRV
XDEC52 WL[105] WL[104] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[5] XPD2[1]
+  S11000X8_XDRV
XDEC53 WL[106] WL[107] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[5] XPD2[1]
+  S11000X8_XDRV
XDEC54 WL[109] WL[108] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[5] XPD2[1]
+  S11000X8_XDRV
XDEC55 WL[110] WL[111] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[5] XPD2[1]
+  S11000X8_XDRV
XDEC56 WL[113] WL[112] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[6] XPD2[1]
+  S11000X8_XDRV
XDEC57 WL[114] WL[115] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[6] XPD2[1]
+  S11000X8_XDRV
XDEC58 WL[117] WL[116] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[6] XPD2[1]
+  S11000X8_XDRV
XDEC59 WL[118] WL[119] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[6] XPD2[1]
+  S11000X8_XDRV
XDEC60 WL[121] WL[120] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[7] XPD2[1]
+  S11000X8_XDRV
XDEC61 WL[122] WL[123] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[7] XPD2[1]
+  S11000X8_XDRV
XDEC62 WL[125] WL[124] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[7] XPD2[1]
+  S11000X8_XDRV
XDEC63 WL[126] WL[127] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[7] XPD2[1]
+  S11000X8_XDRV
XDEC64 WL[129] WL[128] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[2]
+  S11000X8_XDRV
XDEC65 WL[130] WL[131] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[2]
+  S11000X8_XDRV
XDEC66 WL[133] WL[132] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[2]
+  S11000X8_XDRV
XDEC67 WL[134] WL[135] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[2]
+  S11000X8_XDRV
XDEC68 WL[137] WL[136] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[2]
+  S11000X8_XDRV
XDEC69 WL[138] WL[139] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[2]
+  S11000X8_XDRV
XDEC70 WL[141] WL[140] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[2]
+  S11000X8_XDRV
XDEC71 WL[142] WL[143] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[2]
+  S11000X8_XDRV
XDEC72 WL[145] WL[144] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[2]
+  S11000X8_XDRV
XDEC73 WL[146] WL[147] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[2]
+  S11000X8_XDRV
XDEC74 WL[149] WL[148] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[2]
+  S11000X8_XDRV
XDEC75 WL[150] WL[151] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[2]
+  S11000X8_XDRV
XDEC76 WL[153] WL[152] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[2]
+  S11000X8_XDRV
XDEC77 WL[154] WL[155] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[2]
+  S11000X8_XDRV
XDEC78 WL[157] WL[156] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[2]
+  S11000X8_XDRV
XDEC79 WL[158] WL[159] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[2]
+  S11000X8_XDRV
XDEC80 WL[161] WL[160] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[4] XPD2[2]
+  S11000X8_XDRV
XDEC81 WL[162] WL[163] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[4] XPD2[2]
+  S11000X8_XDRV
XDEC82 WL[165] WL[164] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[4] XPD2[2]
+  S11000X8_XDRV
XDEC83 WL[166] WL[167] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[4] XPD2[2]
+  S11000X8_XDRV
XDEC84 WL[169] WL[168] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[5] XPD2[2]
+  S11000X8_XDRV
XDEC85 WL[170] WL[171] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[5] XPD2[2]
+  S11000X8_XDRV
XDEC86 WL[173] WL[172] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[5] XPD2[2]
+  S11000X8_XDRV
XDEC87 WL[174] WL[175] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[5] XPD2[2]
+  S11000X8_XDRV
XDEC88 WL[177] WL[176] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[6] XPD2[2]
+  S11000X8_XDRV
XDEC89 WL[178] WL[179] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[6] XPD2[2]
+  S11000X8_XDRV
XDEC90 WL[181] WL[180] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[6] XPD2[2]
+  S11000X8_XDRV
XDEC91 WL[182] WL[183] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[6] XPD2[2]
+  S11000X8_XDRV
XDEC92 WL[185] WL[184] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[7] XPD2[2]
+  S11000X8_XDRV
XDEC93 WL[186] WL[187] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[7] XPD2[2]
+  S11000X8_XDRV
XDEC94 WL[189] WL[188] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[7] XPD2[2]
+  S11000X8_XDRV
XDEC95 WL[190] WL[191] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[7] XPD2[2]
+  S11000X8_XDRV
XDEC96 WL[193] WL[192] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[3]
+  S11000X8_XDRV
XDEC97 WL[194] WL[195] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[3]
+  S11000X8_XDRV
XDEC98 WL[197] WL[196] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[3]
+  S11000X8_XDRV
XDEC99 WL[198] WL[199] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[3]
+  S11000X8_XDRV
XDEC100 WL[201] WL[200] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[3]
+  S11000X8_XDRV
XDEC101 WL[202] WL[203] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[3]
+  S11000X8_XDRV
XDEC102 WL[205] WL[204] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[3]
+  S11000X8_XDRV
XDEC103 WL[206] WL[207] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[3]
+  S11000X8_XDRV
XDEC104 WL[209] WL[208] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[3]
+  S11000X8_XDRV
XDEC105 WL[210] WL[211] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[3]
+  S11000X8_XDRV
XDEC106 WL[213] WL[212] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[3]
+  S11000X8_XDRV
XDEC107 WL[214] WL[215] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[3]
+  S11000X8_XDRV
XDEC108 WL[217] WL[216] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[3]
+  S11000X8_XDRV
XDEC109 WL[218] WL[219] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[3]
+  S11000X8_XDRV
XDEC110 WL[221] WL[220] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[3]
+  S11000X8_XDRV
XDEC111 WL[222] WL[223] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[3]
+  S11000X8_XDRV
XDEC112 WL[225] WL[224] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[4] XPD2[3]
+  S11000X8_XDRV
XDEC113 WL[226] WL[227] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[4] XPD2[3]
+  S11000X8_XDRV
XDEC114 WL[229] WL[228] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[4] XPD2[3]
+  S11000X8_XDRV
XDEC115 WL[230] WL[231] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[4] XPD2[3]
+  S11000X8_XDRV
XDEC116 WL[233] WL[232] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[5] XPD2[3]
+  S11000X8_XDRV
XDEC117 WL[234] WL[235] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[5] XPD2[3]
+  S11000X8_XDRV
XDEC118 WL[237] WL[236] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[5] XPD2[3]
+  S11000X8_XDRV
XDEC119 WL[238] WL[239] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[5] XPD2[3]
+  S11000X8_XDRV
XDEC120 WL[241] WL[240] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[6] XPD2[3]
+  S11000X8_XDRV
XDEC121 WL[242] WL[243] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[6] XPD2[3]
+  S11000X8_XDRV
XDEC122 WL[245] WL[244] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[6] XPD2[3]
+  S11000X8_XDRV
XDEC123 WL[246] WL[247] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[6] XPD2[3]
+  S11000X8_XDRV
XDEC124 WL[249] WL[248] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[7] XPD2[3]
+  S11000X8_XDRV
XDEC125 WL[250] WL[251] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[7] XPD2[3]
+  S11000X8_XDRV
XDEC126 WL[253] WL[252] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[7] XPD2[3]
+  S11000X8_XDRV
XDEC127 WL[254] WL[255] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[7] XPD2[3]
+  S11000X8_XDRV
XDEC128 WL[257] WL[256] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[4]
+  S11000X8_XDRV
XDEC129 WL[258] WL[259] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[4]
+  S11000X8_XDRV
XDEC130 WL[261] WL[260] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[4]
+  S11000X8_XDRV
XDEC131 WL[262] WL[263] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[4]
+  S11000X8_XDRV
XDEC132 WL[265] WL[264] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[4]
+  S11000X8_XDRV
XDEC133 WL[266] WL[267] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[4]
+  S11000X8_XDRV
XDEC134 WL[269] WL[268] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[4]
+  S11000X8_XDRV
XDEC135 WL[270] WL[271] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[4]
+  S11000X8_XDRV
XDEC136 WL[273] WL[272] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[4]
+  S11000X8_XDRV
XDEC137 WL[274] WL[275] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[4]
+  S11000X8_XDRV
XDEC138 WL[277] WL[276] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[4]
+  S11000X8_XDRV
XDEC139 WL[278] WL[279] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[4]
+  S11000X8_XDRV
XDEC140 WL[281] WL[280] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[4]
+  S11000X8_XDRV
XDEC141 WL[282] WL[283] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[4]
+  S11000X8_XDRV
XDEC142 WL[285] WL[284] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[4]
+  S11000X8_XDRV
XDEC143 WL[286] WL[287] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[4]
+  S11000X8_XDRV
XDEC144 WL[289] WL[288] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[4] XPD2[4]
+  S11000X8_XDRV
XDEC145 WL[290] WL[291] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[4] XPD2[4]
+  S11000X8_XDRV
XDEC146 WL[293] WL[292] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[4] XPD2[4]
+  S11000X8_XDRV
XDEC147 WL[294] WL[295] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[4] XPD2[4]
+  S11000X8_XDRV
XDEC148 WL[297] WL[296] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[5] XPD2[4]
+  S11000X8_XDRV
XDEC149 WL[298] WL[299] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[5] XPD2[4]
+  S11000X8_XDRV
XDEC150 WL[301] WL[300] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[5] XPD2[4]
+  S11000X8_XDRV
XDEC151 WL[302] WL[303] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[5] XPD2[4]
+  S11000X8_XDRV
XDEC152 WL[305] WL[304] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[6] XPD2[4]
+  S11000X8_XDRV
XDEC153 WL[306] WL[307] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[6] XPD2[4]
+  S11000X8_XDRV
XDEC154 WL[309] WL[308] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[6] XPD2[4]
+  S11000X8_XDRV
XDEC155 WL[310] WL[311] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[6] XPD2[4]
+  S11000X8_XDRV
XDEC156 WL[313] WL[312] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[7] XPD2[4]
+  S11000X8_XDRV
XDEC157 WL[314] WL[315] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[7] XPD2[4]
+  S11000X8_XDRV
XDEC158 WL[317] WL[316] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[7] XPD2[4]
+  S11000X8_XDRV
XDEC159 WL[318] WL[319] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[7] XPD2[4]
+  S11000X8_XDRV
XDEC160 WL[321] WL[320] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[5]
+  S11000X8_XDRV
XDEC161 WL[322] WL[323] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[5]
+  S11000X8_XDRV
XDEC162 WL[325] WL[324] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[5]
+  S11000X8_XDRV
XDEC163 WL[326] WL[327] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[5]
+  S11000X8_XDRV
XDEC164 WL[329] WL[328] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[5]
+  S11000X8_XDRV
XDEC165 WL[330] WL[331] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[5]
+  S11000X8_XDRV
XDEC166 WL[333] WL[332] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[5]
+  S11000X8_XDRV
XDEC167 WL[334] WL[335] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[5]
+  S11000X8_XDRV
XDEC168 WL[337] WL[336] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[5]
+  S11000X8_XDRV
XDEC169 WL[338] WL[339] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[5]
+  S11000X8_XDRV
XDEC170 WL[341] WL[340] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[5]
+  S11000X8_XDRV
XDEC171 WL[342] WL[343] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[5]
+  S11000X8_XDRV
XDEC172 WL[345] WL[344] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[5]
+  S11000X8_XDRV
XDEC173 WL[346] WL[347] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[5]
+  S11000X8_XDRV
XDEC174 WL[349] WL[348] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[5]
+  S11000X8_XDRV
XDEC175 WL[350] WL[351] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[5]
+  S11000X8_XDRV
XDEC176 WL[353] WL[352] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[4] XPD2[5]
+  S11000X8_XDRV
XDEC177 WL[354] WL[355] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[4] XPD2[5]
+  S11000X8_XDRV
XDEC178 WL[357] WL[356] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[4] XPD2[5]
+  S11000X8_XDRV
XDEC179 WL[358] WL[359] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[4] XPD2[5]
+  S11000X8_XDRV
XDEC180 WL[361] WL[360] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[5] XPD2[5]
+  S11000X8_XDRV
XDEC181 WL[362] WL[363] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[5] XPD2[5]
+  S11000X8_XDRV
XDEC182 WL[365] WL[364] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[5] XPD2[5]
+  S11000X8_XDRV
XDEC183 WL[366] WL[367] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[5] XPD2[5]
+  S11000X8_XDRV
XDEC184 WL[369] WL[368] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[6] XPD2[5]
+  S11000X8_XDRV
XDEC185 WL[370] WL[371] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[6] XPD2[5]
+  S11000X8_XDRV
XDEC186 WL[373] WL[372] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[6] XPD2[5]
+  S11000X8_XDRV
XDEC187 WL[374] WL[375] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[6] XPD2[5]
+  S11000X8_XDRV
XDEC188 WL[377] WL[376] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[7] XPD2[5]
+  S11000X8_XDRV
XDEC189 WL[378] WL[379] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[7] XPD2[5]
+  S11000X8_XDRV
XDEC190 WL[381] WL[380] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[7] XPD2[5]
+  S11000X8_XDRV
XDEC191 WL[382] WL[383] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[7] XPD2[5]
+  S11000X8_XDRV
XDEC192 WL[385] WL[384] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[6]
+  S11000X8_XDRV
XDEC193 WL[386] WL[387] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[6]
+  S11000X8_XDRV
XDEC194 WL[389] WL[388] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[6]
+  S11000X8_XDRV
XDEC195 WL[390] WL[391] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[6]
+  S11000X8_XDRV
XDEC196 WL[393] WL[392] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[6]
+  S11000X8_XDRV
XDEC197 WL[394] WL[395] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[6]
+  S11000X8_XDRV
XDEC198 WL[397] WL[396] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[6]
+  S11000X8_XDRV
XDEC199 WL[398] WL[399] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[6]
+  S11000X8_XDRV
XDEC200 WL[401] WL[400] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[6]
+  S11000X8_XDRV
XDEC201 WL[402] WL[403] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[6]
+  S11000X8_XDRV
XDEC202 WL[405] WL[404] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[6]
+  S11000X8_XDRV
XDEC203 WL[406] WL[407] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[6]
+  S11000X8_XDRV
XDEC204 WL[409] WL[408] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[6]
+  S11000X8_XDRV
XDEC205 WL[410] WL[411] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[6]
+  S11000X8_XDRV
XDEC206 WL[413] WL[412] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[6]
+  S11000X8_XDRV
XDEC207 WL[414] WL[415] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[6]
+  S11000X8_XDRV
XDEC208 WL[417] WL[416] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[4] XPD2[6]
+  S11000X8_XDRV
XDEC209 WL[418] WL[419] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[4] XPD2[6]
+  S11000X8_XDRV
XDEC210 WL[421] WL[420] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[4] XPD2[6]
+  S11000X8_XDRV
XDEC211 WL[422] WL[423] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[4] XPD2[6]
+  S11000X8_XDRV
XDEC212 WL[425] WL[424] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[5] XPD2[6]
+  S11000X8_XDRV
XDEC213 WL[426] WL[427] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[5] XPD2[6]
+  S11000X8_XDRV
XDEC214 WL[429] WL[428] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[5] XPD2[6]
+  S11000X8_XDRV
XDEC215 WL[430] WL[431] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[5] XPD2[6]
+  S11000X8_XDRV
XDEC216 WL[433] WL[432] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[6] XPD2[6]
+  S11000X8_XDRV
XDEC217 WL[434] WL[435] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[6] XPD2[6]
+  S11000X8_XDRV
XDEC218 WL[437] WL[436] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[6] XPD2[6]
+  S11000X8_XDRV
XDEC219 WL[438] WL[439] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[6] XPD2[6]
+  S11000X8_XDRV
XDEC220 WL[441] WL[440] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[7] XPD2[6]
+  S11000X8_XDRV
XDEC221 WL[442] WL[443] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[7] XPD2[6]
+  S11000X8_XDRV
XDEC222 WL[445] WL[444] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[7] XPD2[6]
+  S11000X8_XDRV
XDEC223 WL[446] WL[447] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[7] XPD2[6]
+  S11000X8_XDRV
XDEC224 WL[449] WL[448] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[0] XPD2[7]
+  S11000X8_XDRV
XDEC225 WL[450] WL[451] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[0] XPD2[7]
+  S11000X8_XDRV
XDEC226 WL[453] WL[452] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[0] XPD2[7]
+  S11000X8_XDRV
XDEC227 WL[454] WL[455] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[0] XPD2[7]
+  S11000X8_XDRV
XDEC228 WL[457] WL[456] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[1] XPD2[7]
+  S11000X8_XDRV
XDEC229 WL[458] WL[459] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[1] XPD2[7]
+  S11000X8_XDRV
XDEC230 WL[461] WL[460] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[1] XPD2[7]
+  S11000X8_XDRV
XDEC231 WL[462] WL[463] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[1] XPD2[7]
+  S11000X8_XDRV
XDEC232 WL[465] WL[464] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[2] XPD2[7]
+  S11000X8_XDRV
XDEC233 WL[466] WL[467] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[2] XPD2[7]
+  S11000X8_XDRV
XDEC234 WL[469] WL[468] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[2] XPD2[7]
+  S11000X8_XDRV
XDEC235 WL[470] WL[471] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[2] XPD2[7]
+  S11000X8_XDRV
XDEC236 WL[473] WL[472] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[3] XPD2[7]
+  S11000X8_XDRV
XDEC237 WL[474] WL[475] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[3] XPD2[7]
+  S11000X8_XDRV
XDEC238 WL[477] WL[476] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[3] XPD2[7]
+  S11000X8_XDRV
XDEC239 WL[478] WL[479] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[3] XPD2[7]
+  S11000X8_XDRV
XDEC240 WL[481] WL[480] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[4] XPD2[7]
+  S11000X8_XDRV
XDEC241 WL[482] WL[483] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[4] XPD2[7]
+  S11000X8_XDRV
XDEC242 WL[485] WL[484] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[4] XPD2[7]
+  S11000X8_XDRV
XDEC243 WL[486] WL[487] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[4] XPD2[7]
+  S11000X8_XDRV
XDEC244 WL[489] WL[488] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[5] XPD2[7]
+  S11000X8_XDRV
XDEC245 WL[490] WL[491] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[5] XPD2[7]
+  S11000X8_XDRV
XDEC246 WL[493] WL[492] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[5] XPD2[7]
+  S11000X8_XDRV
XDEC247 WL[494] WL[495] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[5] XPD2[7]
+  S11000X8_XDRV
XDEC248 WL[497] WL[496] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[6] XPD2[7]
+  S11000X8_XDRV
XDEC249 WL[498] WL[499] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[6] XPD2[7]
+  S11000X8_XDRV
XDEC250 WL[501] WL[500] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[6] XPD2[7]
+  S11000X8_XDRV
XDEC251 WL[502] WL[503] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[6] XPD2[7]
+  S11000X8_XDRV
XDEC252 WL[505] WL[504] WLPY WLPYB0 WLPYB1 XPD0[0] XPD0[1] XPD1[7] XPD2[7]
+  S11000X8_XDRV
XDEC253 WL[506] WL[507] WLPY WLPYB0 WLPYB1 XPD0[3] XPD0[2] XPD1[7] XPD2[7]
+  S11000X8_XDRV
XDEC254 WL[509] WL[508] WLPY WLPYB0 WLPYB1 XPD0[4] XPD0[5] XPD1[7] XPD2[7]
+  S11000X8_XDRV
XDEC255 WL[510] WL[511] WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD1[7] XPD2[7]
+  S11000X8_XDRV
.ENDS

.SUBCKT S11000X8_TRKCOL TRKBL TIEL TRKBLB TRKWL WL[511] WL[510] WL[509] 
+ WL[508] WL[507] WL[506] WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] 
+ WL[499] WL[498] WL[497] WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] 
+ WL[490] WL[489] WL[488] WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] 
+ WL[481] WL[480] WL[479] WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] 
+ WL[472] WL[471] WL[470] WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] 
+ WL[463] WL[462] WL[461] WL[460] WL[459] WL[458] WL[457] WL[456] WL[455] 
+ WL[454] WL[453] WL[452] WL[451] WL[450] WL[449] WL[448] WL[447] WL[446] 
+ WL[445] WL[444] WL[443] WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] 
+ WL[436] WL[435] WL[434] WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] 
+ WL[427] WL[426] WL[425] WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] 
+ WL[418] WL[417] WL[416] WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] 
+ WL[409] WL[408] WL[407] WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] 
+ WL[400] WL[399] WL[398] WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] 
+ WL[391] WL[390] WL[389] WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] 
+ WL[382] WL[381] WL[380] WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] 
+ WL[373] WL[372] WL[371] WL[370] WL[369] WL[368] WL[367] WL[366] WL[365] 
+ WL[364] WL[363] WL[362] WL[361] WL[360] WL[359] WL[358] WL[357] WL[356] 
+ WL[355] WL[354] WL[353] WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] 
+ WL[346] WL[345] WL[344] WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] 
+ WL[337] WL[336] WL[335] WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] 
+ WL[328] WL[327] WL[326] WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] 
+ WL[319] WL[318] WL[317] WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] 
+ WL[310] WL[309] WL[308] WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] 
+ WL[301] WL[300] WL[299] WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] 
+ WL[292] WL[291] WL[290] WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] 
+ WL[283] WL[282] WL[281] WL[280] WL[279] WL[278] WL[277] WL[276] WL[275] 
+ WL[274] WL[273] WL[272] WL[271] WL[270] WL[269] WL[268] WL[267] WL[266] 
+ WL[265] WL[264] WL[263] WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] 
+ WL[256] WL[255] WL[254] WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] 
+ WL[247] WL[246] WL[245] WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] 
+ WL[238] WL[237] WL[236] WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] 
+ WL[229] WL[228] WL[227] WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] 
+ WL[220] WL[219] WL[218] WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] 
+ WL[211] WL[210] WL[209] WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] 
+ WL[202] WL[201] WL[200] WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] 
+ WL[193] WL[192] WL[191] WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] 
+ WL[184] WL[183] WL[182] WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] 
+ WL[175] WL[174] WL[173] WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] 
+ WL[166] WL[165] WL[164] WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] 
+ WL[157] WL[156] WL[155] WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] 
+ WL[148] WL[147] WL[146] WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] 
+ WL[139] WL[138] WL[137] WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] 
+ WL[130] WL[129] WL[128] WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] 
+ WL[121] WL[120] WL[119] WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] 
+ WL[112] WL[111] WL[110] WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] 
+ WL[103] WL[102] WL[101] WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] 
+ WL[93] WL[92] WL[91] WL[90] WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] 
+ WL[82] WL[81] WL[80] WL[79] WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] 
+ WL[71] WL[70] WL[69] WL[68] WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] 
+ WL[60] WL[59] WL[58] WL[57] WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] 
+ WL[49] WL[48] WL[47] WL[46] WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] 
+ WL[38] WL[37] WL[36] WL[35] WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] 
+ WL[27] WL[26] WL[25] WL[24] WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] 
+ WL[16] WL[15] WL[14] WL[13] WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] 
+ WL[5] WL[4] WL[3] WL[2] WL[1] WL[0]
XTRKDUM0 EDG32[1] EDG32[2] TRKBL TIEL WL[1] WL[0] S11000X8_TRKDUMX2
XTRKDUM2 EDG32[2] EDG32[3] TRKBL TIEL WL[3] WL[2] S11000X8_TRKDUMX2
XTRKDUM4 EDG32[3] EDG32[4] TRKBL TIEL WL[5] WL[4] S11000X8_TRKDUMX2
XTRKDUM6 EDG32[4] EDG32[5] TRKBL TIEL WL[7] WL[6] S11000X8_TRKDUMX2
XTRKDUM8 EDG32[5] EDG32[6] TRKBL TIEL WL[9] WL[8] S11000X8_TRKDUMX2
XTRKDUM10 EDG32[6] EDG32[7] TRKBL TIEL WL[11] WL[10] S11000X8_TRKDUMX2
XTRKDUM12 EDG32[7] EDG32[8] TRKBL TIEL WL[13] WL[12] S11000X8_TRKDUMX2
XTRKDUM14 EDG32[8] EDG32[9] TRKBL TIEL WL[15] WL[14] S11000X8_TRKDUMX2
XTRKDUM16 EDG32[9] EDG32[10] TRKBL TIEL WL[17] WL[16] S11000X8_TRKDUMX2
XTRKDUM18 EDG32[10] EDG32[11] TRKBL TIEL WL[19] WL[18] S11000X8_TRKDUMX2
XTRKDUM20 EDG32[11] EDG32[12] TRKBL TIEL WL[21] WL[20] S11000X8_TRKDUMX2
XTRKDUM22 EDG32[12] EDG32[13] TRKBL TIEL WL[23] WL[22] S11000X8_TRKDUMX2
XTRKDUM24 EDG32[13] EDG32[14] TRKBL TIEL WL[25] WL[24] S11000X8_TRKDUMX2
XTRKDUM26 EDG32[14] EDG32[15] TRKBL TIEL WL[27] WL[26] S11000X8_TRKDUMX2
XTRKDUM28 EDG32[15] EDG32[16] TRKBL TIEL WL[29] WL[28] S11000X8_TRKDUMX2
XTRKDUM30 EDG32[16] EDG32[17] TRKBL TIEL WL[31] WL[30] S11000X8_TRKDUMX2
XTRKDUM32 EDG32[17] EDG32[18] TRKBL TIEL WL[33] WL[32] S11000X8_TRKDUMX2
XTRKDUM34 EDG32[18] EDG32[19] TRKBL TIEL WL[35] WL[34] S11000X8_TRKDUMX2
XTRKDUM36 EDG32[19] EDG32[20] TRKBL TIEL WL[37] WL[36] S11000X8_TRKDUMX2
XTRKDUM38 EDG32[20] EDG32[21] TRKBL TIEL WL[39] WL[38] S11000X8_TRKDUMX2
XTRKDUM40 EDG32[21] EDG32[22] TRKBL TIEL WL[41] WL[40] S11000X8_TRKDUMX2
XTRKDUM42 EDG32[22] EDG32[23] TRKBL TIEL WL[43] WL[42] S11000X8_TRKDUMX2
XTRKDUM44 EDG32[23] EDG32[24] TRKBL TIEL WL[45] WL[44] S11000X8_TRKDUMX2
XTRKDUM46 EDG32[24] EDG32[25] TRKBL TIEL WL[47] WL[46] S11000X8_TRKDUMX2
XTRKDUM48 EDG32[25] EDG32[26] TRKBL TIEL WL[49] WL[48] S11000X8_TRKDUMX2
XTRKDUM50 EDG32[26] EDG32[27] TRKBL TIEL WL[51] WL[50] S11000X8_TRKDUMX2
XTRKDUM52 EDG32[27] EDG32[28] TRKBL TIEL WL[53] WL[52] S11000X8_TRKDUMX2
XTRKDUM54 EDG32[28] EDG32[29] TRKBL TIEL WL[55] WL[54] S11000X8_TRKDUMX2
XTRKDUM56 EDG32[29] EDG32[30] TRKBL TIEL WL[57] WL[56] S11000X8_TRKDUMX2
XTRKDUM58 EDG32[30] EDG32[31] TRKBL TIEL WL[59] WL[58] S11000X8_TRKDUMX2
XTRKDUM60 EDG32[31] EDG32[32] TRKBL TIEL WL[61] WL[60] S11000X8_TRKDUMX2
XTRKDUM62 EDG32[32] EDG32[33] TRKBL TIEL WL[63] WL[62] S11000X8_TRKDUMX2
XTRKDUM64 EDG32[34] EDG32[35] TRKBL TIEL WL[65] WL[64] S11000X8_TRKDUMX2
XTRKDUM66 EDG32[35] EDG32[36] TRKBL TIEL WL[67] WL[66] S11000X8_TRKDUMX2
XTRKDUM68 EDG32[36] EDG32[37] TRKBL TIEL WL[69] WL[68] S11000X8_TRKDUMX2
XTRKDUM70 EDG32[37] EDG32[38] TRKBL TIEL WL[71] WL[70] S11000X8_TRKDUMX2
XTRKDUM72 EDG32[38] EDG32[39] TRKBL TIEL WL[73] WL[72] S11000X8_TRKDUMX2
XTRKDUM74 EDG32[39] EDG32[40] TRKBL TIEL WL[75] WL[74] S11000X8_TRKDUMX2
XTRKDUM76 EDG32[40] EDG32[41] TRKBL TIEL WL[77] WL[76] S11000X8_TRKDUMX2
XTRKDUM78 EDG32[41] EDG32[42] TRKBL TIEL WL[79] WL[78] S11000X8_TRKDUMX2
XTRKDUM80 EDG32[42] EDG32[43] TRKBL TIEL WL[81] WL[80] S11000X8_TRKDUMX2
XTRKDUM82 EDG32[43] EDG32[44] TRKBL TIEL WL[83] WL[82] S11000X8_TRKDUMX2
XTRKDUM84 EDG32[44] EDG32[45] TRKBL TIEL WL[85] WL[84] S11000X8_TRKDUMX2
XTRKDUM86 EDG32[45] EDG32[46] TRKBL TIEL WL[87] WL[86] S11000X8_TRKDUMX2
XTRKDUM88 EDG32[46] EDG32[47] TRKBL TIEL WL[89] WL[88] S11000X8_TRKDUMX2
XTRKDUM90 EDG32[47] EDG32[48] TRKBL TIEL WL[91] WL[90] S11000X8_TRKDUMX2
XTRKDUM92 EDG32[48] EDG32[49] TRKBL TIEL WL[93] WL[92] S11000X8_TRKDUMX2
XTRKDUM94 EDG32[49] EDG32[50] TRKBL TIEL WL[95] WL[94] S11000X8_TRKDUMX2
XTRKDUM96 EDG32[50] EDG32[51] TRKBL TIEL WL[97] WL[96] S11000X8_TRKDUMX2
XTRKDUM98 EDG32[51] EDG32[52] TRKBL TIEL WL[99] WL[98] S11000X8_TRKDUMX2
XTRKDUM100 EDG32[52] EDG32[53] TRKBL TIEL WL[101] WL[100] S11000X8_TRKDUMX2
XTRKDUM102 EDG32[53] EDG32[54] TRKBL TIEL WL[103] WL[102] S11000X8_TRKDUMX2
XTRKDUM104 EDG32[54] EDG32[55] TRKBL TIEL WL[105] WL[104] S11000X8_TRKDUMX2
XTRKDUM106 EDG32[55] EDG32[56] TRKBL TIEL WL[107] WL[106] S11000X8_TRKDUMX2
XTRKDUM108 EDG32[56] EDG32[57] TRKBL TIEL WL[109] WL[108] S11000X8_TRKDUMX2
XTRKDUM110 EDG32[57] EDG32[58] TRKBL TIEL WL[111] WL[110] S11000X8_TRKDUMX2
XTRKDUM112 EDG32[58] EDG32[59] TRKBL TIEL WL[113] WL[112] S11000X8_TRKDUMX2
XTRKDUM114 EDG32[59] EDG32[60] TRKBL TIEL WL[115] WL[114] S11000X8_TRKDUMX2
XTRKDUM116 EDG32[60] EDG32[61] TRKBL TIEL WL[117] WL[116] S11000X8_TRKDUMX2
XTRKDUM118 EDG32[61] EDG32[62] TRKBL TIEL WL[119] WL[118] S11000X8_TRKDUMX2
XTRKDUM120 EDG32[62] EDG32[63] TRKBL TIEL WL[121] WL[120] S11000X8_TRKDUMX2
XTRKDUM122 EDG32[63] EDG32[64] TRKBL TIEL WL[123] WL[122] S11000X8_TRKDUMX2
XTRKDUM124 EDG32[64] EDG32[65] TRKBL TIEL WL[125] WL[124] S11000X8_TRKDUMX2
XTRKDUM126 EDG32[65] EDG32[66] TRKBL TIEL WL[127] WL[126] S11000X8_TRKDUMX2
XTRKDUM128 EDG32[67] EDG32[68] TRKBL TIEL WL[129] WL[128] S11000X8_TRKDUMX2
XTRKDUM130 EDG32[68] EDG32[69] TRKBL TIEL WL[131] WL[130] S11000X8_TRKDUMX2
XTRKDUM132 EDG32[69] EDG32[70] TRKBL TIEL WL[133] WL[132] S11000X8_TRKDUMX2
XTRKDUM134 EDG32[70] EDG32[71] TRKBL TIEL WL[135] WL[134] S11000X8_TRKDUMX2
XTRKDUM136 EDG32[71] EDG32[72] TRKBL TIEL WL[137] WL[136] S11000X8_TRKDUMX2
XTRKDUM138 EDG32[72] EDG32[73] TRKBL TIEL WL[139] WL[138] S11000X8_TRKDUMX2
XTRKDUM140 EDG32[73] EDG32[74] TRKBL TIEL WL[141] WL[140] S11000X8_TRKDUMX2
XTRKDUM142 EDG32[74] EDG32[75] TRKBL TIEL WL[143] WL[142] S11000X8_TRKDUMX2
XTRKDUM144 EDG32[75] EDG32[76] TRKBL TIEL WL[145] WL[144] S11000X8_TRKDUMX2
XTRKDUM146 EDG32[76] EDG32[77] TRKBL TIEL WL[147] WL[146] S11000X8_TRKDUMX2
XTRKDUM148 EDG32[77] EDG32[78] TRKBL TIEL WL[149] WL[148] S11000X8_TRKDUMX2
XTRKDUM150 EDG32[78] EDG32[79] TRKBL TIEL WL[151] WL[150] S11000X8_TRKDUMX2
XTRKDUM152 EDG32[79] EDG32[80] TRKBL TIEL WL[153] WL[152] S11000X8_TRKDUMX2
XTRKDUM154 EDG32[80] EDG32[81] TRKBL TIEL WL[155] WL[154] S11000X8_TRKDUMX2
XTRKDUM156 EDG32[81] EDG32[82] TRKBL TIEL WL[157] WL[156] S11000X8_TRKDUMX2
XTRKDUM158 EDG32[82] EDG32[83] TRKBL TIEL WL[159] WL[158] S11000X8_TRKDUMX2
XTRKDUM160 EDG32[83] EDG32[84] TRKBL TIEL WL[161] WL[160] S11000X8_TRKDUMX2
XTRKDUM162 EDG32[84] EDG32[85] TRKBL TIEL WL[163] WL[162] S11000X8_TRKDUMX2
XTRKDUM164 EDG32[85] EDG32[86] TRKBL TIEL WL[165] WL[164] S11000X8_TRKDUMX2
XTRKDUM166 EDG32[86] EDG32[87] TRKBL TIEL WL[167] WL[166] S11000X8_TRKDUMX2
XTRKDUM168 EDG32[87] EDG32[88] TRKBL TIEL WL[169] WL[168] S11000X8_TRKDUMX2
XTRKDUM170 EDG32[88] EDG32[89] TRKBL TIEL WL[171] WL[170] S11000X8_TRKDUMX2
XTRKDUM172 EDG32[89] EDG32[90] TRKBL TIEL WL[173] WL[172] S11000X8_TRKDUMX2
XTRKDUM174 EDG32[90] EDG32[91] TRKBL TIEL WL[175] WL[174] S11000X8_TRKDUMX2
XTRKDUM176 EDG32[91] EDG32[92] TRKBL TIEL WL[177] WL[176] S11000X8_TRKDUMX2
XTRKDUM178 EDG32[92] EDG32[93] TRKBL TIEL WL[179] WL[178] S11000X8_TRKDUMX2
XTRKDUM180 EDG32[93] EDG32[94] TRKBL TIEL WL[181] WL[180] S11000X8_TRKDUMX2
XTRKDUM182 EDG32[94] EDG32[95] TRKBL TIEL WL[183] WL[182] S11000X8_TRKDUMX2
XTRKDUM184 EDG32[95] EDG32[96] TRKBL TIEL WL[185] WL[184] S11000X8_TRKDUMX2
XTRKDUM186 EDG32[96] EDG32[97] TRKBL TIEL WL[187] WL[186] S11000X8_TRKDUMX2
XTRKDUM188 EDG32[97] EDG32[98] TRKBL TIEL WL[189] WL[188] S11000X8_TRKDUMX2
XTRKDUM190 EDG32[98] EDG32[99] TRKBL TIEL WL[191] WL[190] S11000X8_TRKDUMX2
XTRKDUM192 EDG32[100] EDG32[101] TRKBL TIEL WL[193] WL[192] S11000X8_TRKDUMX2
XTRKDUM194 EDG32[101] EDG32[102] TRKBL TIEL WL[195] WL[194] S11000X8_TRKDUMX2
XTRKDUM196 EDG32[102] EDG32[103] TRKBL TIEL WL[197] WL[196] S11000X8_TRKDUMX2
XTRKDUM198 EDG32[103] EDG32[104] TRKBL TIEL WL[199] WL[198] S11000X8_TRKDUMX2
XTRKDUM200 EDG32[104] EDG32[105] TRKBL TIEL WL[201] WL[200] S11000X8_TRKDUMX2
XTRKDUM202 EDG32[105] EDG32[106] TRKBL TIEL WL[203] WL[202] S11000X8_TRKDUMX2
XTRKDUM204 EDG32[106] EDG32[107] TRKBL TIEL WL[205] WL[204] S11000X8_TRKDUMX2
XTRKDUM206 EDG32[107] EDG32[108] TRKBL TIEL WL[207] WL[206] S11000X8_TRKDUMX2
XTRKDUM208 EDG32[108] EDG32[109] TRKBL TIEL WL[209] WL[208] S11000X8_TRKDUMX2
XTRKDUM210 EDG32[109] EDG32[110] TRKBL TIEL WL[211] WL[210] S11000X8_TRKDUMX2
XTRKDUM212 EDG32[110] EDG32[111] TRKBL TIEL WL[213] WL[212] S11000X8_TRKDUMX2
XTRKDUM214 EDG32[111] EDG32[112] TRKBL TIEL WL[215] WL[214] S11000X8_TRKDUMX2
XTRKDUM216 EDG32[112] EDG32[113] TRKBL TIEL WL[217] WL[216] S11000X8_TRKDUMX2
XTRKDUM218 EDG32[113] EDG32[114] TRKBL TIEL WL[219] WL[218] S11000X8_TRKDUMX2
XTRKDUM220 EDG32[114] EDG32[115] TRKBL TIEL WL[221] WL[220] S11000X8_TRKDUMX2
XTRKDUM222 EDG32[115] EDG32[116] TRKBL TIEL WL[223] WL[222] S11000X8_TRKDUMX2
XTRKDUM224 EDG32[116] EDG32[117] TRKBL TIEL WL[225] WL[224] S11000X8_TRKDUMX2
XTRKDUM226 EDG32[117] EDG32[118] TRKBL TIEL WL[227] WL[226] S11000X8_TRKDUMX2
XTRKDUM228 EDG32[118] EDG32[119] TRKBL TIEL WL[229] WL[228] S11000X8_TRKDUMX2
XTRKDUM230 EDG32[119] EDG32[120] TRKBL TIEL WL[231] WL[230] S11000X8_TRKDUMX2
XTRKDUM232 EDG32[120] EDG32[121] TRKBL TIEL WL[233] WL[232] S11000X8_TRKDUMX2
XTRKDUM234 EDG32[121] EDG32[122] TRKBL TIEL WL[235] WL[234] S11000X8_TRKDUMX2
XTRKDUM236 EDG32[122] EDG32[123] TRKBL TIEL WL[237] WL[236] S11000X8_TRKDUMX2
XTRKDUM238 EDG32[123] EDG32[124] TRKBL TIEL WL[239] WL[238] S11000X8_TRKDUMX2
XTRKDUM240 EDG32[124] EDG32[125] TRKBL TIEL WL[241] WL[240] S11000X8_TRKDUMX2
XTRKDUM242 EDG32[125] EDG32[126] TRKBL TIEL WL[243] WL[242] S11000X8_TRKDUMX2
XTRKDUM244 EDG32[126] EDG32[127] TRKBL TIEL WL[245] WL[244] S11000X8_TRKDUMX2
XTRKDUM246 EDG32[127] EDG32[128] TRKBL TIEL WL[247] WL[246] S11000X8_TRKDUMX2
XTRKDUM248 EDG32[128] EDG32[129] TRKBL TIEL WL[249] WL[248] S11000X8_TRKDUMX2
XTRKDUM250 EDG32[129] EDG32[130] TRKBL TIEL WL[251] WL[250] S11000X8_TRKDUMX2
XTRKDUM252 EDG32[130] EDG32[131] TRKBL TIEL WL[253] WL[252] S11000X8_TRKDUMX2
XTRKDUM254 EDG32[131] EDG32[132] TRKBL TIEL WL[255] WL[254] S11000X8_TRKDUMX2
XTRKDUM256 EDG32[133] EDG32[134] TRKBL TIEL WL[257] WL[256] S11000X8_TRKDUMX2
XTRKDUM258 EDG32[134] EDG32[135] TRKBL TIEL WL[259] WL[258] S11000X8_TRKDUMX2
XTRKDUM260 EDG32[135] EDG32[136] TRKBL TIEL WL[261] WL[260] S11000X8_TRKDUMX2
XTRKDUM262 EDG32[136] EDG32[137] TRKBL TIEL WL[263] WL[262] S11000X8_TRKDUMX2
XTRKDUM264 EDG32[137] EDG32[138] TRKBL TIEL WL[265] WL[264] S11000X8_TRKDUMX2
XTRKDUM266 EDG32[138] EDG32[139] TRKBL TIEL WL[267] WL[266] S11000X8_TRKDUMX2
XTRKDUM268 EDG32[139] EDG32[140] TRKBL TIEL WL[269] WL[268] S11000X8_TRKDUMX2
XTRKDUM270 EDG32[140] EDG32[141] TRKBL TIEL WL[271] WL[270] S11000X8_TRKDUMX2
XTRKDUM272 EDG32[141] EDG32[142] TRKBL TIEL WL[273] WL[272] S11000X8_TRKDUMX2
XTRKDUM274 EDG32[142] EDG32[143] TRKBL TIEL WL[275] WL[274] S11000X8_TRKDUMX2
XTRKDUM276 EDG32[143] EDG32[144] TRKBL TIEL WL[277] WL[276] S11000X8_TRKDUMX2
XTRKDUM278 EDG32[144] EDG32[145] TRKBL TIEL WL[279] WL[278] S11000X8_TRKDUMX2
XTRKDUM280 EDG32[145] EDG32[146] TRKBL TIEL WL[281] WL[280] S11000X8_TRKDUMX2
XTRKDUM282 EDG32[146] EDG32[147] TRKBL TIEL WL[283] WL[282] S11000X8_TRKDUMX2
XTRKDUM284 EDG32[147] EDG32[148] TRKBL TIEL WL[285] WL[284] S11000X8_TRKDUMX2
XTRKDUM286 EDG32[148] EDG32[149] TRKBL TIEL WL[287] WL[286] S11000X8_TRKDUMX2
XTRKDUM288 EDG32[149] EDG32[150] TRKBL TIEL WL[289] WL[288] S11000X8_TRKDUMX2
XTRKDUM290 EDG32[150] EDG32[151] TRKBL TIEL WL[291] WL[290] S11000X8_TRKDUMX2
XTRKDUM292 EDG32[151] EDG32[152] TRKBL TIEL WL[293] WL[292] S11000X8_TRKDUMX2
XTRKDUM294 EDG32[152] EDG32[153] TRKBL TIEL WL[295] WL[294] S11000X8_TRKDUMX2
XTRKDUM296 EDG32[153] EDG32[154] TRKBL TIEL WL[297] WL[296] S11000X8_TRKDUMX2
XTRKDUM298 EDG32[154] EDG32[155] TRKBL TIEL WL[299] WL[298] S11000X8_TRKDUMX2
XTRKDUM300 EDG32[155] EDG32[156] TRKBL TIEL WL[301] WL[300] S11000X8_TRKDUMX2
XTRKDUM302 EDG32[156] EDG32[157] TRKBL TIEL WL[303] WL[302] S11000X8_TRKDUMX2
XTRKDUM304 EDG32[157] EDG32[158] TRKBL TIEL WL[305] WL[304] S11000X8_TRKDUMX2
XTRKDUM306 EDG32[158] EDG32[159] TRKBL TIEL WL[307] WL[306] S11000X8_TRKDUMX2
XTRKDUM308 EDG32[159] EDG32[160] TRKBL TIEL WL[309] WL[308] S11000X8_TRKDUMX2
XTRKDUM310 EDG32[160] EDG32[161] TRKBL TIEL WL[311] WL[310] S11000X8_TRKDUMX2
XTRKDUM312 EDG32[161] EDG32[162] TRKBL TIEL WL[313] WL[312] S11000X8_TRKDUMX2
XTRKDUM314 EDG32[162] EDG32[163] TRKBL TIEL WL[315] WL[314] S11000X8_TRKDUMX2
XTRKDUM316 EDG32[163] EDG32[164] TRKBL TIEL WL[317] WL[316] S11000X8_TRKDUMX2
XTRKDUM318 EDG32[164] EDG32[165] TRKBL TIEL WL[319] WL[318] S11000X8_TRKDUMX2
XTRKDUM320 EDG32[166] EDG32[167] TRKBL TIEL WL[321] WL[320] S11000X8_TRKDUMX2
XTRKDUM322 EDG32[167] EDG32[168] TRKBL TIEL WL[323] WL[322] S11000X8_TRKDUMX2
XTRKDUM324 EDG32[168] EDG32[169] TRKBL TIEL WL[325] WL[324] S11000X8_TRKDUMX2
XTRKDUM326 EDG32[169] EDG32[170] TRKBL TIEL WL[327] WL[326] S11000X8_TRKDUMX2
XTRKDUM328 EDG32[170] EDG32[171] TRKBL TIEL WL[329] WL[328] S11000X8_TRKDUMX2
XTRKDUM330 EDG32[171] EDG32[172] TRKBL TIEL WL[331] WL[330] S11000X8_TRKDUMX2
XTRKDUM332 EDG32[172] EDG32[173] TRKBL TIEL WL[333] WL[332] S11000X8_TRKDUMX2
XTRKDUM334 EDG32[173] EDG32[174] TRKBL TIEL WL[335] WL[334] S11000X8_TRKDUMX2
XTRKDUM336 EDG32[174] EDG32[175] TRKBL TIEL WL[337] WL[336] S11000X8_TRKDUMX2
XTRKDUM338 EDG32[175] EDG32[176] TRKBL TIEL WL[339] WL[338] S11000X8_TRKDUMX2
XTRKDUM340 EDG32[176] EDG32[177] TRKBL TIEL WL[341] WL[340] S11000X8_TRKDUMX2
XTRKDUM342 EDG32[177] EDG32[178] TRKBL TIEL WL[343] WL[342] S11000X8_TRKDUMX2
XTRKDUM344 EDG32[178] EDG32[179] TRKBL TIEL WL[345] WL[344] S11000X8_TRKDUMX2
XTRKDUM346 EDG32[179] EDG32[180] TRKBL TIEL WL[347] WL[346] S11000X8_TRKDUMX2
XTRKDUM348 EDG32[180] EDG32[181] TRKBL TIEL WL[349] WL[348] S11000X8_TRKDUMX2
XTRKDUM350 EDG32[181] EDG32[182] TRKBL TIEL WL[351] WL[350] S11000X8_TRKDUMX2
XTRKDUM352 EDG32[182] EDG32[183] TRKBL TIEL WL[353] WL[352] S11000X8_TRKDUMX2
XTRKDUM354 EDG32[183] EDG32[184] TRKBL TIEL WL[355] WL[354] S11000X8_TRKDUMX2
XTRKDUM356 EDG32[184] EDG32[185] TRKBL TIEL WL[357] WL[356] S11000X8_TRKDUMX2
XTRKDUM358 EDG32[185] EDG32[186] TRKBL TIEL WL[359] WL[358] S11000X8_TRKDUMX2
XTRKDUM360 EDG32[186] EDG32[187] TRKBL TIEL WL[361] WL[360] S11000X8_TRKDUMX2
XTRKDUM362 EDG32[187] EDG32[188] TRKBL TIEL WL[363] WL[362] S11000X8_TRKDUMX2
XTRKDUM364 EDG32[188] EDG32[189] TRKBL TIEL WL[365] WL[364] S11000X8_TRKDUMX2
XTRKDUM366 EDG32[189] EDG32[190] TRKBL TIEL WL[367] WL[366] S11000X8_TRKDUMX2
XTRKDUM368 EDG32[190] EDG32[191] TRKBL TIEL WL[369] WL[368] S11000X8_TRKDUMX2
XTRKDUM370 EDG32[191] EDG32[192] TRKBL TIEL WL[371] WL[370] S11000X8_TRKDUMX2
XTRKDUM372 EDG32[192] EDG32[193] TRKBL TIEL WL[373] WL[372] S11000X8_TRKDUMX2
XTRKDUM374 EDG32[193] EDG32[194] TRKBL TIEL WL[375] WL[374] S11000X8_TRKDUMX2
XTRKDUM376 EDG32[194] EDG32[195] TRKBL TIEL WL[377] WL[376] S11000X8_TRKDUMX2
XTRKDUM378 EDG32[195] EDG32[196] TRKBL TIEL WL[379] WL[378] S11000X8_TRKDUMX2
XTRKDUM380 EDG32[196] EDG32[197] TRKBL TIEL WL[381] WL[380] S11000X8_TRKDUMX2
XTRKDUM382 EDG32[197] EDG32[198] TRKBL TIEL WL[383] WL[382] S11000X8_TRKDUMX2
XTRKDUM384 EDG32[199] EDG32[200] TRKBL TIEL WL[385] WL[384] S11000X8_TRKDUMX2
XTRKDUM386 EDG32[200] EDG32[201] TRKBL TIEL WL[387] WL[386] S11000X8_TRKDUMX2
XTRKDUM388 EDG32[201] EDG32[202] TRKBL TIEL WL[389] WL[388] S11000X8_TRKDUMX2
XTRKDUM390 EDG32[202] EDG32[203] TRKBL TIEL WL[391] WL[390] S11000X8_TRKDUMX2
XTRKDUM392 EDG32[203] EDG32[204] TRKBL TIEL WL[393] WL[392] S11000X8_TRKDUMX2
XTRKDUM394 EDG32[204] EDG32[205] TRKBL TIEL WL[395] WL[394] S11000X8_TRKDUMX2
XTRKDUM396 EDG32[205] EDG32[206] TRKBL TIEL WL[397] WL[396] S11000X8_TRKDUMX2
XTRKDUM398 EDG32[206] EDG32[207] TRKBL TIEL WL[399] WL[398] S11000X8_TRKDUMX2
XTRKDUM400 EDG32[207] EDG32[208] TRKBL TIEL WL[401] WL[400] S11000X8_TRKDUMX2
XTRKDUM402 EDG32[208] EDG32[209] TRKBL TIEL WL[403] WL[402] S11000X8_TRKDUMX2
XTRKDUM404 EDG32[209] EDG32[210] TRKBL TIEL WL[405] WL[404] S11000X8_TRKDUMX2
XTRKDUM406 EDG32[210] EDG32[211] TRKBL TIEL WL[407] WL[406] S11000X8_TRKDUMX2
XTRKDUM408 EDG32[211] EDG32[212] TRKBL TIEL WL[409] WL[408] S11000X8_TRKDUMX2
XTRKDUM410 EDG32[212] EDG32[213] TRKBL TIEL WL[411] WL[410] S11000X8_TRKDUMX2
XTRKDUM412 EDG32[213] EDG32[214] TRKBL TIEL WL[413] WL[412] S11000X8_TRKDUMX2
XTRKDUM414 EDG32[214] EDG32[215] TRKBL TIEL WL[415] WL[414] S11000X8_TRKDUMX2
XTRKDUM416 EDG32[215] EDG32[216] TRKBL TIEL WL[417] WL[416] S11000X8_TRKDUMX2
XTRKDUM418 EDG32[216] EDG32[217] TRKBL TIEL WL[419] WL[418] S11000X8_TRKDUMX2
XTRKDUM420 EDG32[217] EDG32[218] TRKBL TIEL WL[421] WL[420] S11000X8_TRKDUMX2
XTRKDUM422 EDG32[218] EDG32[219] TRKBL TIEL WL[423] WL[422] S11000X8_TRKDUMX2
XTRKDUM424 EDG32[219] EDG32[220] TRKBL TIEL WL[425] WL[424] S11000X8_TRKDUMX2
XTRKDUM426 EDG32[220] EDG32[221] TRKBL TIEL WL[427] WL[426] S11000X8_TRKDUMX2
XTRKDUM428 EDG32[221] EDG32[222] TRKBL TIEL WL[429] WL[428] S11000X8_TRKDUMX2
XTRKDUM430 EDG32[222] EDG32[223] TRKBL TIEL WL[431] WL[430] S11000X8_TRKDUMX2
XTRKDUM432 EDG32[223] EDG32[224] TRKBL TIEL WL[433] WL[432] S11000X8_TRKDUMX2
XTRKDUM434 EDG32[224] EDG32[225] TRKBL TIEL WL[435] WL[434] S11000X8_TRKDUMX2
XTRKDUM436 EDG32[225] EDG32[226] TRKBL TIEL WL[437] WL[436] S11000X8_TRKDUMX2
XTRKDUM438 EDG32[226] EDG32[227] TRKBL TIEL WL[439] WL[438] S11000X8_TRKDUMX2
XTRKDUM440 EDG32[227] EDG32[228] TRKBL TIEL WL[441] WL[440] S11000X8_TRKDUMX2
XTRKDUM442 EDG32[228] EDG32[229] TRKBL TIEL WL[443] WL[442] S11000X8_TRKDUMX2
XTRKDUM444 EDG32[229] EDG32[230] TRKBL TIEL WL[445] WL[444] S11000X8_TRKDUMX2
XTRKDUM446 EDG32[230] EDG32[231] TRKBL TIEL WL[447] WL[446] S11000X8_TRKDUMX2
XTRKDUM448 EDG32[232] EDG32[233] TRKBL TIEL WL[449] WL[448] S11000X8_TRKDUMX2
XTRKDUM450 EDG32[233] EDG32[234] TRKBL TIEL WL[451] WL[450] S11000X8_TRKDUMX2
XTRKDUM452 EDG32[234] EDG32[235] TRKBL TIEL WL[453] WL[452] S11000X8_TRKDUMX2
XTRKDUM454 EDG32[235] EDG32[236] TRKBL TIEL WL[455] WL[454] S11000X8_TRKDUMX2
XTRKDUM456 EDG32[236] EDG32[237] TRKBL TIEL WL[457] WL[456] S11000X8_TRKDUMX2
XTRKDUM458 EDG32[237] EDG32[238] TRKBL TIEL WL[459] WL[458] S11000X8_TRKDUMX2
XTRKDUM460 EDG32[238] EDG32[239] TRKBL TIEL WL[461] WL[460] S11000X8_TRKDUMX2
XTRKDUM462 EDG32[239] EDG32[240] TRKBL TIEL WL[463] WL[462] S11000X8_TRKDUMX2
XTRKDUM464 EDG32[240] EDG32[241] TRKBL TIEL WL[465] WL[464] S11000X8_TRKDUMX2
XTRKDUM466 EDG32[241] EDG32[242] TRKBL TIEL WL[467] WL[466] S11000X8_TRKDUMX2
XTRKDUM468 EDG32[242] EDG32[243] TRKBL TIEL WL[469] WL[468] S11000X8_TRKDUMX2
XTRKDUM470 EDG32[243] EDG32[244] TRKBL TIEL WL[471] WL[470] S11000X8_TRKDUMX2
XTRKDUM472 EDG32[244] EDG32[245] TRKBL TIEL WL[473] WL[472] S11000X8_TRKDUMX2
XTRKDUM474 EDG32[245] EDG32[246] TRKBL TIEL WL[475] WL[474] S11000X8_TRKDUMX2
XTRKDUM476 EDG32[246] EDG32[247] TRKBL TIEL WL[477] WL[476] S11000X8_TRKDUMX2
XTRKDUM478 EDG32[247] EDG32[248] TRKBL TIEL WL[479] WL[478] S11000X8_TRKDUMX2
XTRKDUM480 EDG32[248] EDG32[249] TRKBL TIEL WL[481] WL[480] S11000X8_TRKDUMX2
XTRKDUM482 EDG32[249] EDG32[250] TRKBL TIEL WL[483] WL[482] S11000X8_TRKDUMX2
XTRKDUM484 EDG32[250] EDG32[251] TRKBL TIEL WL[485] WL[484] S11000X8_TRKDUMX2
XTRKDUM486 EDG32[251] EDG32[252] TRKBL TIEL WL[487] WL[486] S11000X8_TRKDUMX2
XTRKDUM488 EDG32[252] EDG32[253] TRKBL TIEL WL[489] WL[488] S11000X8_TRKDUMX2
XTRKDUM490 EDG32[253] EDG32[254] TRKBL TIEL WL[491] WL[490] S11000X8_TRKDUMX2
XTRKDUM492 EDG32[254] EDG32[255] TRKBL TIEL WL[493] WL[492] S11000X8_TRKDUMX2
XTRKDUM494 EDG32[255] EDG32[256] TRKBL TIEL WL[495] WL[494] S11000X8_TRKDUMX2
XTRKDUM496 EDG32[256] EDG32[257] TRKBL TIEL WL[497] WL[496] S11000X8_TRKDUMX2
XTRKDUM498 EDG32[257] EDG32[258] TRKBL TIEL WL[499] WL[498] S11000X8_TRKDUMX2
XTRKDUM500 EDG32[258] EDG32[259] TRKBL TIEL WL[501] WL[500] S11000X8_TRKDUMX2
XTRKNOR502 EDG32[259] EDG32[260] TRKBL TRKBLB TRKWL WL[503] WL[502]
+  S11000X8_TRKNORX2
XTRKNOR504 EDG32[260] EDG32[261] TRKBL TRKBLB TRKWL WL[505] WL[504]
+  S11000X8_TRKNORX2
XTRKNOR506 EDG32[261] EDG32[262] TRKBL TRKBLB TRKWL WL[507] WL[506]
+  S11000X8_TRKNORX2
XTRKNOR508 EDG32[262] EDG32[263] TRKBL TRKBLB TRKWL WL[509] WL[508]
+  S11000X8_TRKNORX2
XTRKNOR510 EDG32[263] EDG32[264] TRKBL TRKBLB TRKWL WL[511] WL[510]
+  S11000X8_TRKNORX2
.ENDS

.SUBCKT S11000X8_CORECOLUMN BL0 BL1 BLB0 BLB1 WL[0] WL[1] WL[2] WL[3] WL[4] 
+ WL[5] WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] 
+ WL[16] WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] 
+ WL[27] WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] 
+ WL[38] WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] 
+ WL[49] WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] 
+ WL[60] WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] 
+ WL[71] WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] 
+ WL[82] WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] 
+ WL[93] WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] 
+ WL[103] WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] 
+ WL[112] WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] 
+ WL[121] WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] 
+ WL[130] WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] 
+ WL[139] WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] 
+ WL[148] WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] 
+ WL[157] WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] 
+ WL[166] WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] 
+ WL[175] WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] 
+ WL[184] WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] 
+ WL[193] WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] 
+ WL[202] WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] 
+ WL[211] WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] 
+ WL[220] WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] 
+ WL[229] WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] 
+ WL[238] WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] 
+ WL[247] WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] 
+ WL[256] WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] 
+ WL[265] WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] 
+ WL[274] WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] 
+ WL[283] WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] 
+ WL[292] WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] 
+ WL[301] WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] 
+ WL[310] WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] 
+ WL[319] WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] 
+ WL[328] WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] 
+ WL[337] WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] 
+ WL[346] WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] 
+ WL[355] WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] 
+ WL[364] WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] 
+ WL[373] WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] 
+ WL[382] WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] 
+ WL[391] WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] 
+ WL[400] WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] 
+ WL[409] WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] 
+ WL[418] WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] 
+ WL[427] WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] 
+ WL[436] WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] 
+ WL[445] WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] 
+ WL[454] WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] 
+ WL[463] WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] 
+ WL[472] WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] 
+ WL[481] WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] 
+ WL[490] WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] 
+ WL[499] WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] 
+ WL[508] WL[509] WL[510] WL[511]
XBITCELLX2_0 BL0 BL1 BLB0 BLB1 WL[0] WL[1] S11000X8_CELLX4
XBITCELLX2_1 BL0 BL1 BLB0 BLB1 WL[2] WL[3] S11000X8_CELLX4
XBITCELLX2_2 BL0 BL1 BLB0 BLB1 WL[4] WL[5] S11000X8_CELLX4
XBITCELLX2_3 BL0 BL1 BLB0 BLB1 WL[6] WL[7] S11000X8_CELLX4
XBITCELLX2_4 BL0 BL1 BLB0 BLB1 WL[8] WL[9] S11000X8_CELLX4
XBITCELLX2_5 BL0 BL1 BLB0 BLB1 WL[10] WL[11] S11000X8_CELLX4
XBITCELLX2_6 BL0 BL1 BLB0 BLB1 WL[12] WL[13] S11000X8_CELLX4
XBITCELLX2_7 BL0 BL1 BLB0 BLB1 WL[14] WL[15] S11000X8_CELLX4
XBITCELLX2_8 BL0 BL1 BLB0 BLB1 WL[16] WL[17] S11000X8_CELLX4
XBITCELLX2_9 BL0 BL1 BLB0 BLB1 WL[18] WL[19] S11000X8_CELLX4
XBITCELLX2_10 BL0 BL1 BLB0 BLB1 WL[20] WL[21] S11000X8_CELLX4
XBITCELLX2_11 BL0 BL1 BLB0 BLB1 WL[22] WL[23] S11000X8_CELLX4
XBITCELLX2_12 BL0 BL1 BLB0 BLB1 WL[24] WL[25] S11000X8_CELLX4
XBITCELLX2_13 BL0 BL1 BLB0 BLB1 WL[26] WL[27] S11000X8_CELLX4
XBITCELLX2_14 BL0 BL1 BLB0 BLB1 WL[28] WL[29] S11000X8_CELLX4
XBITCELLX2_15 BL0 BL1 BLB0 BLB1 WL[30] WL[31] S11000X8_CELLX4
XBITCELLX2_16 BL0 BL1 BLB0 BLB1 WL[32] WL[33] S11000X8_CELLX4
XBITCELLX2_17 BL0 BL1 BLB0 BLB1 WL[34] WL[35] S11000X8_CELLX4
XBITCELLX2_18 BL0 BL1 BLB0 BLB1 WL[36] WL[37] S11000X8_CELLX4
XBITCELLX2_19 BL0 BL1 BLB0 BLB1 WL[38] WL[39] S11000X8_CELLX4
XBITCELLX2_20 BL0 BL1 BLB0 BLB1 WL[40] WL[41] S11000X8_CELLX4
XBITCELLX2_21 BL0 BL1 BLB0 BLB1 WL[42] WL[43] S11000X8_CELLX4
XBITCELLX2_22 BL0 BL1 BLB0 BLB1 WL[44] WL[45] S11000X8_CELLX4
XBITCELLX2_23 BL0 BL1 BLB0 BLB1 WL[46] WL[47] S11000X8_CELLX4
XBITCELLX2_24 BL0 BL1 BLB0 BLB1 WL[48] WL[49] S11000X8_CELLX4
XBITCELLX2_25 BL0 BL1 BLB0 BLB1 WL[50] WL[51] S11000X8_CELLX4
XBITCELLX2_26 BL0 BL1 BLB0 BLB1 WL[52] WL[53] S11000X8_CELLX4
XBITCELLX2_27 BL0 BL1 BLB0 BLB1 WL[54] WL[55] S11000X8_CELLX4
XBITCELLX2_28 BL0 BL1 BLB0 BLB1 WL[56] WL[57] S11000X8_CELLX4
XBITCELLX2_29 BL0 BL1 BLB0 BLB1 WL[58] WL[59] S11000X8_CELLX4
XBITCELLX2_30 BL0 BL1 BLB0 BLB1 WL[60] WL[61] S11000X8_CELLX4
XBITCELLX2_31 BL0 BL1 BLB0 BLB1 WL[62] WL[63] S11000X8_CELLX4
XBITCELLX2_32 BL0 BL1 BLB0 BLB1 WL[64] WL[65] S11000X8_CELLX4
XBITCELLX2_33 BL0 BL1 BLB0 BLB1 WL[66] WL[67] S11000X8_CELLX4
XBITCELLX2_34 BL0 BL1 BLB0 BLB1 WL[68] WL[69] S11000X8_CELLX4
XBITCELLX2_35 BL0 BL1 BLB0 BLB1 WL[70] WL[71] S11000X8_CELLX4
XBITCELLX2_36 BL0 BL1 BLB0 BLB1 WL[72] WL[73] S11000X8_CELLX4
XBITCELLX2_37 BL0 BL1 BLB0 BLB1 WL[74] WL[75] S11000X8_CELLX4
XBITCELLX2_38 BL0 BL1 BLB0 BLB1 WL[76] WL[77] S11000X8_CELLX4
XBITCELLX2_39 BL0 BL1 BLB0 BLB1 WL[78] WL[79] S11000X8_CELLX4
XBITCELLX2_40 BL0 BL1 BLB0 BLB1 WL[80] WL[81] S11000X8_CELLX4
XBITCELLX2_41 BL0 BL1 BLB0 BLB1 WL[82] WL[83] S11000X8_CELLX4
XBITCELLX2_42 BL0 BL1 BLB0 BLB1 WL[84] WL[85] S11000X8_CELLX4
XBITCELLX2_43 BL0 BL1 BLB0 BLB1 WL[86] WL[87] S11000X8_CELLX4
XBITCELLX2_44 BL0 BL1 BLB0 BLB1 WL[88] WL[89] S11000X8_CELLX4
XBITCELLX2_45 BL0 BL1 BLB0 BLB1 WL[90] WL[91] S11000X8_CELLX4
XBITCELLX2_46 BL0 BL1 BLB0 BLB1 WL[92] WL[93] S11000X8_CELLX4
XBITCELLX2_47 BL0 BL1 BLB0 BLB1 WL[94] WL[95] S11000X8_CELLX4
XBITCELLX2_48 BL0 BL1 BLB0 BLB1 WL[96] WL[97] S11000X8_CELLX4
XBITCELLX2_49 BL0 BL1 BLB0 BLB1 WL[98] WL[99] S11000X8_CELLX4
XBITCELLX2_50 BL0 BL1 BLB0 BLB1 WL[100] WL[101] S11000X8_CELLX4
XBITCELLX2_51 BL0 BL1 BLB0 BLB1 WL[102] WL[103] S11000X8_CELLX4
XBITCELLX2_52 BL0 BL1 BLB0 BLB1 WL[104] WL[105] S11000X8_CELLX4
XBITCELLX2_53 BL0 BL1 BLB0 BLB1 WL[106] WL[107] S11000X8_CELLX4
XBITCELLX2_54 BL0 BL1 BLB0 BLB1 WL[108] WL[109] S11000X8_CELLX4
XBITCELLX2_55 BL0 BL1 BLB0 BLB1 WL[110] WL[111] S11000X8_CELLX4
XBITCELLX2_56 BL0 BL1 BLB0 BLB1 WL[112] WL[113] S11000X8_CELLX4
XBITCELLX2_57 BL0 BL1 BLB0 BLB1 WL[114] WL[115] S11000X8_CELLX4
XBITCELLX2_58 BL0 BL1 BLB0 BLB1 WL[116] WL[117] S11000X8_CELLX4
XBITCELLX2_59 BL0 BL1 BLB0 BLB1 WL[118] WL[119] S11000X8_CELLX4
XBITCELLX2_60 BL0 BL1 BLB0 BLB1 WL[120] WL[121] S11000X8_CELLX4
XBITCELLX2_61 BL0 BL1 BLB0 BLB1 WL[122] WL[123] S11000X8_CELLX4
XBITCELLX2_62 BL0 BL1 BLB0 BLB1 WL[124] WL[125] S11000X8_CELLX4
XBITCELLX2_63 BL0 BL1 BLB0 BLB1 WL[126] WL[127] S11000X8_CELLX4
XBITCELLX2_64 BL0 BL1 BLB0 BLB1 WL[128] WL[129] S11000X8_CELLX4
XBITCELLX2_65 BL0 BL1 BLB0 BLB1 WL[130] WL[131] S11000X8_CELLX4
XBITCELLX2_66 BL0 BL1 BLB0 BLB1 WL[132] WL[133] S11000X8_CELLX4
XBITCELLX2_67 BL0 BL1 BLB0 BLB1 WL[134] WL[135] S11000X8_CELLX4
XBITCELLX2_68 BL0 BL1 BLB0 BLB1 WL[136] WL[137] S11000X8_CELLX4
XBITCELLX2_69 BL0 BL1 BLB0 BLB1 WL[138] WL[139] S11000X8_CELLX4
XBITCELLX2_70 BL0 BL1 BLB0 BLB1 WL[140] WL[141] S11000X8_CELLX4
XBITCELLX2_71 BL0 BL1 BLB0 BLB1 WL[142] WL[143] S11000X8_CELLX4
XBITCELLX2_72 BL0 BL1 BLB0 BLB1 WL[144] WL[145] S11000X8_CELLX4
XBITCELLX2_73 BL0 BL1 BLB0 BLB1 WL[146] WL[147] S11000X8_CELLX4
XBITCELLX2_74 BL0 BL1 BLB0 BLB1 WL[148] WL[149] S11000X8_CELLX4
XBITCELLX2_75 BL0 BL1 BLB0 BLB1 WL[150] WL[151] S11000X8_CELLX4
XBITCELLX2_76 BL0 BL1 BLB0 BLB1 WL[152] WL[153] S11000X8_CELLX4
XBITCELLX2_77 BL0 BL1 BLB0 BLB1 WL[154] WL[155] S11000X8_CELLX4
XBITCELLX2_78 BL0 BL1 BLB0 BLB1 WL[156] WL[157] S11000X8_CELLX4
XBITCELLX2_79 BL0 BL1 BLB0 BLB1 WL[158] WL[159] S11000X8_CELLX4
XBITCELLX2_80 BL0 BL1 BLB0 BLB1 WL[160] WL[161] S11000X8_CELLX4
XBITCELLX2_81 BL0 BL1 BLB0 BLB1 WL[162] WL[163] S11000X8_CELLX4
XBITCELLX2_82 BL0 BL1 BLB0 BLB1 WL[164] WL[165] S11000X8_CELLX4
XBITCELLX2_83 BL0 BL1 BLB0 BLB1 WL[166] WL[167] S11000X8_CELLX4
XBITCELLX2_84 BL0 BL1 BLB0 BLB1 WL[168] WL[169] S11000X8_CELLX4
XBITCELLX2_85 BL0 BL1 BLB0 BLB1 WL[170] WL[171] S11000X8_CELLX4
XBITCELLX2_86 BL0 BL1 BLB0 BLB1 WL[172] WL[173] S11000X8_CELLX4
XBITCELLX2_87 BL0 BL1 BLB0 BLB1 WL[174] WL[175] S11000X8_CELLX4
XBITCELLX2_88 BL0 BL1 BLB0 BLB1 WL[176] WL[177] S11000X8_CELLX4
XBITCELLX2_89 BL0 BL1 BLB0 BLB1 WL[178] WL[179] S11000X8_CELLX4
XBITCELLX2_90 BL0 BL1 BLB0 BLB1 WL[180] WL[181] S11000X8_CELLX4
XBITCELLX2_91 BL0 BL1 BLB0 BLB1 WL[182] WL[183] S11000X8_CELLX4
XBITCELLX2_92 BL0 BL1 BLB0 BLB1 WL[184] WL[185] S11000X8_CELLX4
XBITCELLX2_93 BL0 BL1 BLB0 BLB1 WL[186] WL[187] S11000X8_CELLX4
XBITCELLX2_94 BL0 BL1 BLB0 BLB1 WL[188] WL[189] S11000X8_CELLX4
XBITCELLX2_95 BL0 BL1 BLB0 BLB1 WL[190] WL[191] S11000X8_CELLX4
XBITCELLX2_96 BL0 BL1 BLB0 BLB1 WL[192] WL[193] S11000X8_CELLX4
XBITCELLX2_97 BL0 BL1 BLB0 BLB1 WL[194] WL[195] S11000X8_CELLX4
XBITCELLX2_98 BL0 BL1 BLB0 BLB1 WL[196] WL[197] S11000X8_CELLX4
XBITCELLX2_99 BL0 BL1 BLB0 BLB1 WL[198] WL[199] S11000X8_CELLX4
XBITCELLX2_100 BL0 BL1 BLB0 BLB1 WL[200] WL[201] S11000X8_CELLX4
XBITCELLX2_101 BL0 BL1 BLB0 BLB1 WL[202] WL[203] S11000X8_CELLX4
XBITCELLX2_102 BL0 BL1 BLB0 BLB1 WL[204] WL[205] S11000X8_CELLX4
XBITCELLX2_103 BL0 BL1 BLB0 BLB1 WL[206] WL[207] S11000X8_CELLX4
XBITCELLX2_104 BL0 BL1 BLB0 BLB1 WL[208] WL[209] S11000X8_CELLX4
XBITCELLX2_105 BL0 BL1 BLB0 BLB1 WL[210] WL[211] S11000X8_CELLX4
XBITCELLX2_106 BL0 BL1 BLB0 BLB1 WL[212] WL[213] S11000X8_CELLX4
XBITCELLX2_107 BL0 BL1 BLB0 BLB1 WL[214] WL[215] S11000X8_CELLX4
XBITCELLX2_108 BL0 BL1 BLB0 BLB1 WL[216] WL[217] S11000X8_CELLX4
XBITCELLX2_109 BL0 BL1 BLB0 BLB1 WL[218] WL[219] S11000X8_CELLX4
XBITCELLX2_110 BL0 BL1 BLB0 BLB1 WL[220] WL[221] S11000X8_CELLX4
XBITCELLX2_111 BL0 BL1 BLB0 BLB1 WL[222] WL[223] S11000X8_CELLX4
XBITCELLX2_112 BL0 BL1 BLB0 BLB1 WL[224] WL[225] S11000X8_CELLX4
XBITCELLX2_113 BL0 BL1 BLB0 BLB1 WL[226] WL[227] S11000X8_CELLX4
XBITCELLX2_114 BL0 BL1 BLB0 BLB1 WL[228] WL[229] S11000X8_CELLX4
XBITCELLX2_115 BL0 BL1 BLB0 BLB1 WL[230] WL[231] S11000X8_CELLX4
XBITCELLX2_116 BL0 BL1 BLB0 BLB1 WL[232] WL[233] S11000X8_CELLX4
XBITCELLX2_117 BL0 BL1 BLB0 BLB1 WL[234] WL[235] S11000X8_CELLX4
XBITCELLX2_118 BL0 BL1 BLB0 BLB1 WL[236] WL[237] S11000X8_CELLX4
XBITCELLX2_119 BL0 BL1 BLB0 BLB1 WL[238] WL[239] S11000X8_CELLX4
XBITCELLX2_120 BL0 BL1 BLB0 BLB1 WL[240] WL[241] S11000X8_CELLX4
XBITCELLX2_121 BL0 BL1 BLB0 BLB1 WL[242] WL[243] S11000X8_CELLX4
XBITCELLX2_122 BL0 BL1 BLB0 BLB1 WL[244] WL[245] S11000X8_CELLX4
XBITCELLX2_123 BL0 BL1 BLB0 BLB1 WL[246] WL[247] S11000X8_CELLX4
XBITCELLX2_124 BL0 BL1 BLB0 BLB1 WL[248] WL[249] S11000X8_CELLX4
XBITCELLX2_125 BL0 BL1 BLB0 BLB1 WL[250] WL[251] S11000X8_CELLX4
XBITCELLX2_126 BL0 BL1 BLB0 BLB1 WL[252] WL[253] S11000X8_CELLX4
XBITCELLX2_127 BL0 BL1 BLB0 BLB1 WL[254] WL[255] S11000X8_CELLX4
XBITCELLX2_128 BL0 BL1 BLB0 BLB1 WL[256] WL[257] S11000X8_CELLX4
XBITCELLX2_129 BL0 BL1 BLB0 BLB1 WL[258] WL[259] S11000X8_CELLX4
XBITCELLX2_130 BL0 BL1 BLB0 BLB1 WL[260] WL[261] S11000X8_CELLX4
XBITCELLX2_131 BL0 BL1 BLB0 BLB1 WL[262] WL[263] S11000X8_CELLX4
XBITCELLX2_132 BL0 BL1 BLB0 BLB1 WL[264] WL[265] S11000X8_CELLX4
XBITCELLX2_133 BL0 BL1 BLB0 BLB1 WL[266] WL[267] S11000X8_CELLX4
XBITCELLX2_134 BL0 BL1 BLB0 BLB1 WL[268] WL[269] S11000X8_CELLX4
XBITCELLX2_135 BL0 BL1 BLB0 BLB1 WL[270] WL[271] S11000X8_CELLX4
XBITCELLX2_136 BL0 BL1 BLB0 BLB1 WL[272] WL[273] S11000X8_CELLX4
XBITCELLX2_137 BL0 BL1 BLB0 BLB1 WL[274] WL[275] S11000X8_CELLX4
XBITCELLX2_138 BL0 BL1 BLB0 BLB1 WL[276] WL[277] S11000X8_CELLX4
XBITCELLX2_139 BL0 BL1 BLB0 BLB1 WL[278] WL[279] S11000X8_CELLX4
XBITCELLX2_140 BL0 BL1 BLB0 BLB1 WL[280] WL[281] S11000X8_CELLX4
XBITCELLX2_141 BL0 BL1 BLB0 BLB1 WL[282] WL[283] S11000X8_CELLX4
XBITCELLX2_142 BL0 BL1 BLB0 BLB1 WL[284] WL[285] S11000X8_CELLX4
XBITCELLX2_143 BL0 BL1 BLB0 BLB1 WL[286] WL[287] S11000X8_CELLX4
XBITCELLX2_144 BL0 BL1 BLB0 BLB1 WL[288] WL[289] S11000X8_CELLX4
XBITCELLX2_145 BL0 BL1 BLB0 BLB1 WL[290] WL[291] S11000X8_CELLX4
XBITCELLX2_146 BL0 BL1 BLB0 BLB1 WL[292] WL[293] S11000X8_CELLX4
XBITCELLX2_147 BL0 BL1 BLB0 BLB1 WL[294] WL[295] S11000X8_CELLX4
XBITCELLX2_148 BL0 BL1 BLB0 BLB1 WL[296] WL[297] S11000X8_CELLX4
XBITCELLX2_149 BL0 BL1 BLB0 BLB1 WL[298] WL[299] S11000X8_CELLX4
XBITCELLX2_150 BL0 BL1 BLB0 BLB1 WL[300] WL[301] S11000X8_CELLX4
XBITCELLX2_151 BL0 BL1 BLB0 BLB1 WL[302] WL[303] S11000X8_CELLX4
XBITCELLX2_152 BL0 BL1 BLB0 BLB1 WL[304] WL[305] S11000X8_CELLX4
XBITCELLX2_153 BL0 BL1 BLB0 BLB1 WL[306] WL[307] S11000X8_CELLX4
XBITCELLX2_154 BL0 BL1 BLB0 BLB1 WL[308] WL[309] S11000X8_CELLX4
XBITCELLX2_155 BL0 BL1 BLB0 BLB1 WL[310] WL[311] S11000X8_CELLX4
XBITCELLX2_156 BL0 BL1 BLB0 BLB1 WL[312] WL[313] S11000X8_CELLX4
XBITCELLX2_157 BL0 BL1 BLB0 BLB1 WL[314] WL[315] S11000X8_CELLX4
XBITCELLX2_158 BL0 BL1 BLB0 BLB1 WL[316] WL[317] S11000X8_CELLX4
XBITCELLX2_159 BL0 BL1 BLB0 BLB1 WL[318] WL[319] S11000X8_CELLX4
XBITCELLX2_160 BL0 BL1 BLB0 BLB1 WL[320] WL[321] S11000X8_CELLX4
XBITCELLX2_161 BL0 BL1 BLB0 BLB1 WL[322] WL[323] S11000X8_CELLX4
XBITCELLX2_162 BL0 BL1 BLB0 BLB1 WL[324] WL[325] S11000X8_CELLX4
XBITCELLX2_163 BL0 BL1 BLB0 BLB1 WL[326] WL[327] S11000X8_CELLX4
XBITCELLX2_164 BL0 BL1 BLB0 BLB1 WL[328] WL[329] S11000X8_CELLX4
XBITCELLX2_165 BL0 BL1 BLB0 BLB1 WL[330] WL[331] S11000X8_CELLX4
XBITCELLX2_166 BL0 BL1 BLB0 BLB1 WL[332] WL[333] S11000X8_CELLX4
XBITCELLX2_167 BL0 BL1 BLB0 BLB1 WL[334] WL[335] S11000X8_CELLX4
XBITCELLX2_168 BL0 BL1 BLB0 BLB1 WL[336] WL[337] S11000X8_CELLX4
XBITCELLX2_169 BL0 BL1 BLB0 BLB1 WL[338] WL[339] S11000X8_CELLX4
XBITCELLX2_170 BL0 BL1 BLB0 BLB1 WL[340] WL[341] S11000X8_CELLX4
XBITCELLX2_171 BL0 BL1 BLB0 BLB1 WL[342] WL[343] S11000X8_CELLX4
XBITCELLX2_172 BL0 BL1 BLB0 BLB1 WL[344] WL[345] S11000X8_CELLX4
XBITCELLX2_173 BL0 BL1 BLB0 BLB1 WL[346] WL[347] S11000X8_CELLX4
XBITCELLX2_174 BL0 BL1 BLB0 BLB1 WL[348] WL[349] S11000X8_CELLX4
XBITCELLX2_175 BL0 BL1 BLB0 BLB1 WL[350] WL[351] S11000X8_CELLX4
XBITCELLX2_176 BL0 BL1 BLB0 BLB1 WL[352] WL[353] S11000X8_CELLX4
XBITCELLX2_177 BL0 BL1 BLB0 BLB1 WL[354] WL[355] S11000X8_CELLX4
XBITCELLX2_178 BL0 BL1 BLB0 BLB1 WL[356] WL[357] S11000X8_CELLX4
XBITCELLX2_179 BL0 BL1 BLB0 BLB1 WL[358] WL[359] S11000X8_CELLX4
XBITCELLX2_180 BL0 BL1 BLB0 BLB1 WL[360] WL[361] S11000X8_CELLX4
XBITCELLX2_181 BL0 BL1 BLB0 BLB1 WL[362] WL[363] S11000X8_CELLX4
XBITCELLX2_182 BL0 BL1 BLB0 BLB1 WL[364] WL[365] S11000X8_CELLX4
XBITCELLX2_183 BL0 BL1 BLB0 BLB1 WL[366] WL[367] S11000X8_CELLX4
XBITCELLX2_184 BL0 BL1 BLB0 BLB1 WL[368] WL[369] S11000X8_CELLX4
XBITCELLX2_185 BL0 BL1 BLB0 BLB1 WL[370] WL[371] S11000X8_CELLX4
XBITCELLX2_186 BL0 BL1 BLB0 BLB1 WL[372] WL[373] S11000X8_CELLX4
XBITCELLX2_187 BL0 BL1 BLB0 BLB1 WL[374] WL[375] S11000X8_CELLX4
XBITCELLX2_188 BL0 BL1 BLB0 BLB1 WL[376] WL[377] S11000X8_CELLX4
XBITCELLX2_189 BL0 BL1 BLB0 BLB1 WL[378] WL[379] S11000X8_CELLX4
XBITCELLX2_190 BL0 BL1 BLB0 BLB1 WL[380] WL[381] S11000X8_CELLX4
XBITCELLX2_191 BL0 BL1 BLB0 BLB1 WL[382] WL[383] S11000X8_CELLX4
XBITCELLX2_192 BL0 BL1 BLB0 BLB1 WL[384] WL[385] S11000X8_CELLX4
XBITCELLX2_193 BL0 BL1 BLB0 BLB1 WL[386] WL[387] S11000X8_CELLX4
XBITCELLX2_194 BL0 BL1 BLB0 BLB1 WL[388] WL[389] S11000X8_CELLX4
XBITCELLX2_195 BL0 BL1 BLB0 BLB1 WL[390] WL[391] S11000X8_CELLX4
XBITCELLX2_196 BL0 BL1 BLB0 BLB1 WL[392] WL[393] S11000X8_CELLX4
XBITCELLX2_197 BL0 BL1 BLB0 BLB1 WL[394] WL[395] S11000X8_CELLX4
XBITCELLX2_198 BL0 BL1 BLB0 BLB1 WL[396] WL[397] S11000X8_CELLX4
XBITCELLX2_199 BL0 BL1 BLB0 BLB1 WL[398] WL[399] S11000X8_CELLX4
XBITCELLX2_200 BL0 BL1 BLB0 BLB1 WL[400] WL[401] S11000X8_CELLX4
XBITCELLX2_201 BL0 BL1 BLB0 BLB1 WL[402] WL[403] S11000X8_CELLX4
XBITCELLX2_202 BL0 BL1 BLB0 BLB1 WL[404] WL[405] S11000X8_CELLX4
XBITCELLX2_203 BL0 BL1 BLB0 BLB1 WL[406] WL[407] S11000X8_CELLX4
XBITCELLX2_204 BL0 BL1 BLB0 BLB1 WL[408] WL[409] S11000X8_CELLX4
XBITCELLX2_205 BL0 BL1 BLB0 BLB1 WL[410] WL[411] S11000X8_CELLX4
XBITCELLX2_206 BL0 BL1 BLB0 BLB1 WL[412] WL[413] S11000X8_CELLX4
XBITCELLX2_207 BL0 BL1 BLB0 BLB1 WL[414] WL[415] S11000X8_CELLX4
XBITCELLX2_208 BL0 BL1 BLB0 BLB1 WL[416] WL[417] S11000X8_CELLX4
XBITCELLX2_209 BL0 BL1 BLB0 BLB1 WL[418] WL[419] S11000X8_CELLX4
XBITCELLX2_210 BL0 BL1 BLB0 BLB1 WL[420] WL[421] S11000X8_CELLX4
XBITCELLX2_211 BL0 BL1 BLB0 BLB1 WL[422] WL[423] S11000X8_CELLX4
XBITCELLX2_212 BL0 BL1 BLB0 BLB1 WL[424] WL[425] S11000X8_CELLX4
XBITCELLX2_213 BL0 BL1 BLB0 BLB1 WL[426] WL[427] S11000X8_CELLX4
XBITCELLX2_214 BL0 BL1 BLB0 BLB1 WL[428] WL[429] S11000X8_CELLX4
XBITCELLX2_215 BL0 BL1 BLB0 BLB1 WL[430] WL[431] S11000X8_CELLX4
XBITCELLX2_216 BL0 BL1 BLB0 BLB1 WL[432] WL[433] S11000X8_CELLX4
XBITCELLX2_217 BL0 BL1 BLB0 BLB1 WL[434] WL[435] S11000X8_CELLX4
XBITCELLX2_218 BL0 BL1 BLB0 BLB1 WL[436] WL[437] S11000X8_CELLX4
XBITCELLX2_219 BL0 BL1 BLB0 BLB1 WL[438] WL[439] S11000X8_CELLX4
XBITCELLX2_220 BL0 BL1 BLB0 BLB1 WL[440] WL[441] S11000X8_CELLX4
XBITCELLX2_221 BL0 BL1 BLB0 BLB1 WL[442] WL[443] S11000X8_CELLX4
XBITCELLX2_222 BL0 BL1 BLB0 BLB1 WL[444] WL[445] S11000X8_CELLX4
XBITCELLX2_223 BL0 BL1 BLB0 BLB1 WL[446] WL[447] S11000X8_CELLX4
XBITCELLX2_224 BL0 BL1 BLB0 BLB1 WL[448] WL[449] S11000X8_CELLX4
XBITCELLX2_225 BL0 BL1 BLB0 BLB1 WL[450] WL[451] S11000X8_CELLX4
XBITCELLX2_226 BL0 BL1 BLB0 BLB1 WL[452] WL[453] S11000X8_CELLX4
XBITCELLX2_227 BL0 BL1 BLB0 BLB1 WL[454] WL[455] S11000X8_CELLX4
XBITCELLX2_228 BL0 BL1 BLB0 BLB1 WL[456] WL[457] S11000X8_CELLX4
XBITCELLX2_229 BL0 BL1 BLB0 BLB1 WL[458] WL[459] S11000X8_CELLX4
XBITCELLX2_230 BL0 BL1 BLB0 BLB1 WL[460] WL[461] S11000X8_CELLX4
XBITCELLX2_231 BL0 BL1 BLB0 BLB1 WL[462] WL[463] S11000X8_CELLX4
XBITCELLX2_232 BL0 BL1 BLB0 BLB1 WL[464] WL[465] S11000X8_CELLX4
XBITCELLX2_233 BL0 BL1 BLB0 BLB1 WL[466] WL[467] S11000X8_CELLX4
XBITCELLX2_234 BL0 BL1 BLB0 BLB1 WL[468] WL[469] S11000X8_CELLX4
XBITCELLX2_235 BL0 BL1 BLB0 BLB1 WL[470] WL[471] S11000X8_CELLX4
XBITCELLX2_236 BL0 BL1 BLB0 BLB1 WL[472] WL[473] S11000X8_CELLX4
XBITCELLX2_237 BL0 BL1 BLB0 BLB1 WL[474] WL[475] S11000X8_CELLX4
XBITCELLX2_238 BL0 BL1 BLB0 BLB1 WL[476] WL[477] S11000X8_CELLX4
XBITCELLX2_239 BL0 BL1 BLB0 BLB1 WL[478] WL[479] S11000X8_CELLX4
XBITCELLX2_240 BL0 BL1 BLB0 BLB1 WL[480] WL[481] S11000X8_CELLX4
XBITCELLX2_241 BL0 BL1 BLB0 BLB1 WL[482] WL[483] S11000X8_CELLX4
XBITCELLX2_242 BL0 BL1 BLB0 BLB1 WL[484] WL[485] S11000X8_CELLX4
XBITCELLX2_243 BL0 BL1 BLB0 BLB1 WL[486] WL[487] S11000X8_CELLX4
XBITCELLX2_244 BL0 BL1 BLB0 BLB1 WL[488] WL[489] S11000X8_CELLX4
XBITCELLX2_245 BL0 BL1 BLB0 BLB1 WL[490] WL[491] S11000X8_CELLX4
XBITCELLX2_246 BL0 BL1 BLB0 BLB1 WL[492] WL[493] S11000X8_CELLX4
XBITCELLX2_247 BL0 BL1 BLB0 BLB1 WL[494] WL[495] S11000X8_CELLX4
XBITCELLX2_248 BL0 BL1 BLB0 BLB1 WL[496] WL[497] S11000X8_CELLX4
XBITCELLX2_249 BL0 BL1 BLB0 BLB1 WL[498] WL[499] S11000X8_CELLX4
XBITCELLX2_250 BL0 BL1 BLB0 BLB1 WL[500] WL[501] S11000X8_CELLX4
XBITCELLX2_251 BL0 BL1 BLB0 BLB1 WL[502] WL[503] S11000X8_CELLX4
XBITCELLX2_252 BL0 BL1 BLB0 BLB1 WL[504] WL[505] S11000X8_CELLX4
XBITCELLX2_253 BL0 BL1 BLB0 BLB1 WL[506] WL[507] S11000X8_CELLX4
XBITCELLX2_254 BL0 BL1 BLB0 BLB1 WL[508] WL[509] S11000X8_CELLX4
XBITCELLX2_255 BL0 BL1 BLB0 BLB1 WL[510] WL[511] S11000X8_CELLX4
.ENDS

.SUBCKT TS1N65LPA4096X8M8 Q[0] Q[1] Q[2] Q[3] Q[4] Q[5] Q[6] Q[7] A[0] A[1] 
+ A[2] A[3] A[4] A[5] A[6] A[7] A[8] A[9] A[10] A[11] BWEB[0] BWEB[1] BWEB[2] 
+ BWEB[3] BWEB[4] BWEB[5] BWEB[6] BWEB[7] CEB CLK D[0] D[1] D[2] D[3] D[4] D[5] 
+ D[6] D[7] WEB TSEL[0] TSEL[1]
XLCOLUMN0 BL[0] BL[1] BLB[0] BLB[1] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] 
+ WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] 
+ WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] 
+ WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] 
+ WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] 
+ WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] 
+ WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] 
+ WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] 
+ WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] 
+ WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] 
+ WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] 
+ WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] 
+ WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] 
+ WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] 
+ WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] 
+ WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] 
+ WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] 
+ WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] 
+ WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] 
+ WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] 
+ WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] 
+ WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] 
+ WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] 
+ WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] 
+ WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] 
+ WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] 
+ WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] 
+ WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] 
+ WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] 
+ WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] 
+ WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] 
+ WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] 
+ WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] 
+ WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] 
+ WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] WL[383] 
+ WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] WL[392] 
+ WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] WL[401] 
+ WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] WL[410] 
+ WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] WL[419] 
+ WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] WL[428] 
+ WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] WL[437] 
+ WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] WL[446] 
+ WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] WL[455] 
+ WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] WL[464] 
+ WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] WL[473] 
+ WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] WL[482] 
+ WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] WL[491] 
+ WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] WL[500] 
+ WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] WL[509] 
+ WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN1 BL[2] BL[3] BLB[2] BLB[3] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] 
+ WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] 
+ WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] 
+ WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] 
+ WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] 
+ WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] 
+ WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] 
+ WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] 
+ WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] 
+ WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] 
+ WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] 
+ WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] 
+ WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] 
+ WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] 
+ WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] 
+ WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] 
+ WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] 
+ WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] 
+ WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] 
+ WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] 
+ WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] 
+ WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] 
+ WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] 
+ WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] 
+ WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] 
+ WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] 
+ WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] 
+ WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] 
+ WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] 
+ WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] 
+ WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] 
+ WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] 
+ WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] 
+ WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] 
+ WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] WL[383] 
+ WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] WL[392] 
+ WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] WL[401] 
+ WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] WL[410] 
+ WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] WL[419] 
+ WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] WL[428] 
+ WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] WL[437] 
+ WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] WL[446] 
+ WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] WL[455] 
+ WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] WL[464] 
+ WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] WL[473] 
+ WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] WL[482] 
+ WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] WL[491] 
+ WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] WL[500] 
+ WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] WL[509] 
+ WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN2 BL[4] BL[5] BLB[4] BLB[5] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] 
+ WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] 
+ WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] 
+ WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] 
+ WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] 
+ WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] 
+ WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] 
+ WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] 
+ WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] 
+ WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] 
+ WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] 
+ WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] 
+ WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] 
+ WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] 
+ WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] 
+ WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] 
+ WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] 
+ WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] 
+ WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] 
+ WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] 
+ WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] 
+ WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] 
+ WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] 
+ WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] 
+ WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] 
+ WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] 
+ WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] 
+ WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] 
+ WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] 
+ WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] 
+ WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] 
+ WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] 
+ WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] 
+ WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] 
+ WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] WL[383] 
+ WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] WL[392] 
+ WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] WL[401] 
+ WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] WL[410] 
+ WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] WL[419] 
+ WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] WL[428] 
+ WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] WL[437] 
+ WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] WL[446] 
+ WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] WL[455] 
+ WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] WL[464] 
+ WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] WL[473] 
+ WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] WL[482] 
+ WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] WL[491] 
+ WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] WL[500] 
+ WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] WL[509] 
+ WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN3 BL[6] BL[7] BLB[6] BLB[7] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] 
+ WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] 
+ WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] 
+ WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] 
+ WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] 
+ WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] 
+ WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] 
+ WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] 
+ WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] 
+ WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] 
+ WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] 
+ WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] 
+ WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] 
+ WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] 
+ WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] 
+ WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] 
+ WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] 
+ WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] 
+ WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] 
+ WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] 
+ WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] 
+ WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] 
+ WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] 
+ WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] 
+ WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] 
+ WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] 
+ WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] 
+ WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] 
+ WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] 
+ WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] 
+ WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] 
+ WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] 
+ WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] 
+ WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] 
+ WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] WL[383] 
+ WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] WL[392] 
+ WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] WL[401] 
+ WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] WL[410] 
+ WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] WL[419] 
+ WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] WL[428] 
+ WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] WL[437] 
+ WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] WL[446] 
+ WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] WL[455] 
+ WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] WL[464] 
+ WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] WL[473] 
+ WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] WL[482] 
+ WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] WL[491] 
+ WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] WL[500] 
+ WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] WL[509] 
+ WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN4 BL[8] BL[9] BLB[8] BLB[9] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] WL[6] 
+ WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] WL[17] 
+ WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] WL[28] 
+ WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] WL[39] 
+ WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] WL[50] 
+ WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] WL[61] 
+ WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] WL[72] 
+ WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] WL[83] 
+ WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] WL[94] 
+ WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] WL[104] 
+ WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] WL[113] 
+ WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] WL[122] 
+ WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] WL[131] 
+ WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] WL[140] 
+ WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] WL[149] 
+ WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] WL[158] 
+ WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] WL[167] 
+ WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] WL[176] 
+ WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] WL[185] 
+ WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] WL[194] 
+ WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] WL[203] 
+ WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] WL[212] 
+ WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] WL[221] 
+ WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] WL[230] 
+ WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] WL[239] 
+ WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] WL[248] 
+ WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] WL[257] 
+ WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] WL[266] 
+ WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] WL[275] 
+ WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] WL[284] 
+ WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] WL[293] 
+ WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] WL[302] 
+ WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] WL[311] 
+ WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] WL[320] 
+ WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] WL[329] 
+ WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] WL[338] 
+ WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] WL[347] 
+ WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] WL[356] 
+ WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] WL[365] 
+ WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] WL[374] 
+ WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] WL[383] 
+ WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] WL[392] 
+ WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] WL[401] 
+ WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] WL[410] 
+ WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] WL[419] 
+ WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] WL[428] 
+ WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] WL[437] 
+ WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] WL[446] 
+ WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] WL[455] 
+ WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] WL[464] 
+ WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] WL[473] 
+ WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] WL[482] 
+ WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] WL[491] 
+ WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] WL[500] 
+ WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] WL[509] 
+ WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN5 BL[10] BL[11] BLB[10] BLB[11] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN6 BL[12] BL[13] BLB[12] BLB[13] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN7 BL[14] BL[15] BLB[14] BLB[15] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN8 BL[16] BL[17] BLB[16] BLB[17] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN9 BL[18] BL[19] BLB[18] BLB[19] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN10 BL[20] BL[21] BLB[20] BLB[21] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN11 BL[22] BL[23] BLB[22] BLB[23] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN12 BL[24] BL[25] BLB[24] BLB[25] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN13 BL[26] BL[27] BLB[26] BLB[27] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN14 BL[28] BL[29] BLB[28] BLB[29] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN15 BL[30] BL[31] BLB[30] BLB[31] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN16 BL[32] BL[33] BLB[32] BLB[33] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN17 BL[34] BL[35] BLB[34] BLB[35] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN18 BL[36] BL[37] BLB[36] BLB[37] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN19 BL[38] BL[39] BLB[38] BLB[39] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN20 BL[40] BL[41] BLB[40] BLB[41] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN21 BL[42] BL[43] BLB[42] BLB[43] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN22 BL[44] BL[45] BLB[44] BLB[45] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN23 BL[46] BL[47] BLB[46] BLB[47] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN24 BL[48] BL[49] BLB[48] BLB[49] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN25 BL[50] BL[51] BLB[50] BLB[51] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN26 BL[52] BL[53] BLB[52] BLB[53] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN27 BL[54] BL[55] BLB[54] BLB[55] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN28 BL[56] BL[57] BLB[56] BLB[57] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN29 BL[58] BL[59] BLB[58] BLB[59] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN30 BL[60] BL[61] BLB[60] BLB[61] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XLCOLUMN31 BL[62] BL[63] BLB[62] BLB[63] WL[0] WL[1] WL[2] WL[3] WL[4] WL[5] 
+ WL[6] WL[7] WL[8] WL[9] WL[10] WL[11] WL[12] WL[13] WL[14] WL[15] WL[16] 
+ WL[17] WL[18] WL[19] WL[20] WL[21] WL[22] WL[23] WL[24] WL[25] WL[26] WL[27] 
+ WL[28] WL[29] WL[30] WL[31] WL[32] WL[33] WL[34] WL[35] WL[36] WL[37] WL[38] 
+ WL[39] WL[40] WL[41] WL[42] WL[43] WL[44] WL[45] WL[46] WL[47] WL[48] WL[49] 
+ WL[50] WL[51] WL[52] WL[53] WL[54] WL[55] WL[56] WL[57] WL[58] WL[59] WL[60] 
+ WL[61] WL[62] WL[63] WL[64] WL[65] WL[66] WL[67] WL[68] WL[69] WL[70] WL[71] 
+ WL[72] WL[73] WL[74] WL[75] WL[76] WL[77] WL[78] WL[79] WL[80] WL[81] WL[82] 
+ WL[83] WL[84] WL[85] WL[86] WL[87] WL[88] WL[89] WL[90] WL[91] WL[92] WL[93] 
+ WL[94] WL[95] WL[96] WL[97] WL[98] WL[99] WL[100] WL[101] WL[102] WL[103] 
+ WL[104] WL[105] WL[106] WL[107] WL[108] WL[109] WL[110] WL[111] WL[112] 
+ WL[113] WL[114] WL[115] WL[116] WL[117] WL[118] WL[119] WL[120] WL[121] 
+ WL[122] WL[123] WL[124] WL[125] WL[126] WL[127] WL[128] WL[129] WL[130] 
+ WL[131] WL[132] WL[133] WL[134] WL[135] WL[136] WL[137] WL[138] WL[139] 
+ WL[140] WL[141] WL[142] WL[143] WL[144] WL[145] WL[146] WL[147] WL[148] 
+ WL[149] WL[150] WL[151] WL[152] WL[153] WL[154] WL[155] WL[156] WL[157] 
+ WL[158] WL[159] WL[160] WL[161] WL[162] WL[163] WL[164] WL[165] WL[166] 
+ WL[167] WL[168] WL[169] WL[170] WL[171] WL[172] WL[173] WL[174] WL[175] 
+ WL[176] WL[177] WL[178] WL[179] WL[180] WL[181] WL[182] WL[183] WL[184] 
+ WL[185] WL[186] WL[187] WL[188] WL[189] WL[190] WL[191] WL[192] WL[193] 
+ WL[194] WL[195] WL[196] WL[197] WL[198] WL[199] WL[200] WL[201] WL[202] 
+ WL[203] WL[204] WL[205] WL[206] WL[207] WL[208] WL[209] WL[210] WL[211] 
+ WL[212] WL[213] WL[214] WL[215] WL[216] WL[217] WL[218] WL[219] WL[220] 
+ WL[221] WL[222] WL[223] WL[224] WL[225] WL[226] WL[227] WL[228] WL[229] 
+ WL[230] WL[231] WL[232] WL[233] WL[234] WL[235] WL[236] WL[237] WL[238] 
+ WL[239] WL[240] WL[241] WL[242] WL[243] WL[244] WL[245] WL[246] WL[247] 
+ WL[248] WL[249] WL[250] WL[251] WL[252] WL[253] WL[254] WL[255] WL[256] 
+ WL[257] WL[258] WL[259] WL[260] WL[261] WL[262] WL[263] WL[264] WL[265] 
+ WL[266] WL[267] WL[268] WL[269] WL[270] WL[271] WL[272] WL[273] WL[274] 
+ WL[275] WL[276] WL[277] WL[278] WL[279] WL[280] WL[281] WL[282] WL[283] 
+ WL[284] WL[285] WL[286] WL[287] WL[288] WL[289] WL[290] WL[291] WL[292] 
+ WL[293] WL[294] WL[295] WL[296] WL[297] WL[298] WL[299] WL[300] WL[301] 
+ WL[302] WL[303] WL[304] WL[305] WL[306] WL[307] WL[308] WL[309] WL[310] 
+ WL[311] WL[312] WL[313] WL[314] WL[315] WL[316] WL[317] WL[318] WL[319] 
+ WL[320] WL[321] WL[322] WL[323] WL[324] WL[325] WL[326] WL[327] WL[328] 
+ WL[329] WL[330] WL[331] WL[332] WL[333] WL[334] WL[335] WL[336] WL[337] 
+ WL[338] WL[339] WL[340] WL[341] WL[342] WL[343] WL[344] WL[345] WL[346] 
+ WL[347] WL[348] WL[349] WL[350] WL[351] WL[352] WL[353] WL[354] WL[355] 
+ WL[356] WL[357] WL[358] WL[359] WL[360] WL[361] WL[362] WL[363] WL[364] 
+ WL[365] WL[366] WL[367] WL[368] WL[369] WL[370] WL[371] WL[372] WL[373] 
+ WL[374] WL[375] WL[376] WL[377] WL[378] WL[379] WL[380] WL[381] WL[382] 
+ WL[383] WL[384] WL[385] WL[386] WL[387] WL[388] WL[389] WL[390] WL[391] 
+ WL[392] WL[393] WL[394] WL[395] WL[396] WL[397] WL[398] WL[399] WL[400] 
+ WL[401] WL[402] WL[403] WL[404] WL[405] WL[406] WL[407] WL[408] WL[409] 
+ WL[410] WL[411] WL[412] WL[413] WL[414] WL[415] WL[416] WL[417] WL[418] 
+ WL[419] WL[420] WL[421] WL[422] WL[423] WL[424] WL[425] WL[426] WL[427] 
+ WL[428] WL[429] WL[430] WL[431] WL[432] WL[433] WL[434] WL[435] WL[436] 
+ WL[437] WL[438] WL[439] WL[440] WL[441] WL[442] WL[443] WL[444] WL[445] 
+ WL[446] WL[447] WL[448] WL[449] WL[450] WL[451] WL[452] WL[453] WL[454] 
+ WL[455] WL[456] WL[457] WL[458] WL[459] WL[460] WL[461] WL[462] WL[463] 
+ WL[464] WL[465] WL[466] WL[467] WL[468] WL[469] WL[470] WL[471] WL[472] 
+ WL[473] WL[474] WL[475] WL[476] WL[477] WL[478] WL[479] WL[480] WL[481] 
+ WL[482] WL[483] WL[484] WL[485] WL[486] WL[487] WL[488] WL[489] WL[490] 
+ WL[491] WL[492] WL[493] WL[494] WL[495] WL[496] WL[497] WL[498] WL[499] 
+ WL[500] WL[501] WL[502] WL[503] WL[504] WL[505] WL[506] WL[507] WL[508] 
+ WL[509] WL[510] WL[511] S11000X8_CORECOLUMN
XIO0 Q[0] BL[0] BL[1] BL[2] BL[3] BL[4] BL[5] BL[6] BL[7] BLB[0] BLB[1] BLB[2] 
+ BLB[3] BLB[4] BLB[5] BLB[6] BLB[7] AWTI BIST_BUF BWEB[0] TIELB D[0] DCLK 
+ TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0] S11000X8_IO_M8
XIO1 Q[1] BL[8] BL[9] BL[10] BL[11] BL[12] BL[13] BL[14] BL[15] BLB[8] BLB[9] 
+ BLB[10] BLB[11] BLB[12] BLB[13] BLB[14] BLB[15] AWTI BIST_BUF BWEB[1] TIELB 
+ D[1] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0]
+  S11000X8_IO_M8
XIO2 Q[2] BL[16] BL[17] BL[18] BL[19] BL[20] BL[21] BL[22] BL[23] BLB[16] 
+ BLB[17] BLB[18] BLB[19] BLB[20] BLB[21] BLB[22] BLB[23] AWTI BIST_BUF BWEB[2]
+ TIELB D[2] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0]
+  S11000X8_IO_M8
XIO3 Q[3] BL[24] BL[25] BL[26] BL[27] BL[28] BL[29] BL[30] BL[31] BLB[24] 
+ BLB[25] BLB[26] BLB[27] BLB[28] BLB[29] BLB[30] BLB[31] AWTI BIST_BUF BWEB[3]
+ TIELB D[3] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0]
+  S11000X8_IO_M8
XIO4 Q[4] BL[32] BL[33] BL[34] BL[35] BL[36] BL[37] BL[38] BL[39] BLB[32] 
+ BLB[33] BLB[34] BLB[35] BLB[36] BLB[37] BLB[38] BLB[39] AWTI BIST_BUF BWEB[4]
+ TIELB D[4] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0]
+  S11000X8_IO_M8
XIO5 Q[5] BL[40] BL[41] BL[42] BL[43] BL[44] BL[45] BL[46] BL[47] BLB[40] 
+ BLB[41] BLB[42] BLB[43] BLB[44] BLB[45] BLB[46] BLB[47] AWTI BIST_BUF BWEB[5]
+ TIELB D[5] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0]
+  S11000X8_IO_M8
XIO6 Q[6] BL[48] BL[49] BL[50] BL[51] BL[52] BL[53] BL[54] BL[55] BLB[48] 
+ BLB[49] BLB[50] BLB[51] BLB[52] BLB[53] BLB[54] BLB[55] AWTI BIST_BUF BWEB[6]
+ TIELB D[6] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0]
+  S11000X8_IO_M8
XIO7 Q[7] BL[56] BL[57] BL[58] BL[59] BL[60] BL[61] BL[62] BL[63] BLB[56] 
+ BLB[57] BLB[58] BLB[59] BLB[60] BLB[61] BLB[62] BLB[63] AWTI BIST_BUF BWEB[7]
+ TIELB D[7] DCLK TIELB GW_RB WLPX Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] Y32[0]
+  S11000X8_IO_M8
XDEC TRKBL TIEH WL[511] WL[510] WL[509] WL[508] WL[507] WL[506] WL[505] 
+ WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] WL[496] 
+ WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] WL[487] 
+ WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] WL[478] 
+ WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] WL[469] 
+ WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] WL[460] 
+ WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] WL[451] 
+ WL[450] WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] WL[442] 
+ WL[441] WL[440] WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] WL[433] 
+ WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426] WL[425] WL[424] 
+ WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416] WL[415] 
+ WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] WL[406] 
+ WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] WL[397] 
+ WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] WL[388] 
+ WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] WL[379] 
+ WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] WL[370] 
+ WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] WL[361] 
+ WL[360] WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] WL[352] 
+ WL[351] WL[350] WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] WL[343] 
+ WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336] WL[335] WL[334] 
+ WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326] WL[325] 
+ WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] WL[316] 
+ WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] WL[307] 
+ WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] WL[298] 
+ WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] WL[289] 
+ WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] WL[280] 
+ WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] WL[271] 
+ WL[270] WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] WL[262] 
+ WL[261] WL[260] WL[259] WL[258] WL[257] WL[256] WL[255] WL[254] WL[253] 
+ WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] WL[244] 
+ WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] WL[235] 
+ WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] WL[226] 
+ WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] WL[217] 
+ WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] WL[208] 
+ WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] WL[199] 
+ WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] WL[190] 
+ WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] WL[181] 
+ WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] WL[172] 
+ WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] WL[163] 
+ WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] WL[154] 
+ WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] WL[145] 
+ WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] WL[136] 
+ WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] WL[127] 
+ WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] WL[118] 
+ WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] WL[109] 
+ WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] WL[100] 
+ WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] WL[89] 
+ WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] WL[78] 
+ WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] WL[67] 
+ WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] WL[56] 
+ WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] WL[45] 
+ WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] WL[34] 
+ WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] WL[23] 
+ WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] WL[12] 
+ WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] WL[0] 
+ TRKWL WLPY WLPYB0 WLPYB1 XPD0[7] XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] 
+ XPD0[1] XPD0[0] XPD1[7] XPD1[6] XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] 
+ XPD1[0] XPD2[7] XPD2[6] XPD2[5] XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0]
+  S11000X8_DECODER
XTRKCOL TRKBL TIEL TIEH TRKWL WL[511] WL[510] WL[509] WL[508] WL[507] WL[506] 
+ WL[505] WL[504] WL[503] WL[502] WL[501] WL[500] WL[499] WL[498] WL[497] 
+ WL[496] WL[495] WL[494] WL[493] WL[492] WL[491] WL[490] WL[489] WL[488] 
+ WL[487] WL[486] WL[485] WL[484] WL[483] WL[482] WL[481] WL[480] WL[479] 
+ WL[478] WL[477] WL[476] WL[475] WL[474] WL[473] WL[472] WL[471] WL[470] 
+ WL[469] WL[468] WL[467] WL[466] WL[465] WL[464] WL[463] WL[462] WL[461] 
+ WL[460] WL[459] WL[458] WL[457] WL[456] WL[455] WL[454] WL[453] WL[452] 
+ WL[451] WL[450] WL[449] WL[448] WL[447] WL[446] WL[445] WL[444] WL[443] 
+ WL[442] WL[441] WL[440] WL[439] WL[438] WL[437] WL[436] WL[435] WL[434] 
+ WL[433] WL[432] WL[431] WL[430] WL[429] WL[428] WL[427] WL[426] WL[425] 
+ WL[424] WL[423] WL[422] WL[421] WL[420] WL[419] WL[418] WL[417] WL[416] 
+ WL[415] WL[414] WL[413] WL[412] WL[411] WL[410] WL[409] WL[408] WL[407] 
+ WL[406] WL[405] WL[404] WL[403] WL[402] WL[401] WL[400] WL[399] WL[398] 
+ WL[397] WL[396] WL[395] WL[394] WL[393] WL[392] WL[391] WL[390] WL[389] 
+ WL[388] WL[387] WL[386] WL[385] WL[384] WL[383] WL[382] WL[381] WL[380] 
+ WL[379] WL[378] WL[377] WL[376] WL[375] WL[374] WL[373] WL[372] WL[371] 
+ WL[370] WL[369] WL[368] WL[367] WL[366] WL[365] WL[364] WL[363] WL[362] 
+ WL[361] WL[360] WL[359] WL[358] WL[357] WL[356] WL[355] WL[354] WL[353] 
+ WL[352] WL[351] WL[350] WL[349] WL[348] WL[347] WL[346] WL[345] WL[344] 
+ WL[343] WL[342] WL[341] WL[340] WL[339] WL[338] WL[337] WL[336] WL[335] 
+ WL[334] WL[333] WL[332] WL[331] WL[330] WL[329] WL[328] WL[327] WL[326] 
+ WL[325] WL[324] WL[323] WL[322] WL[321] WL[320] WL[319] WL[318] WL[317] 
+ WL[316] WL[315] WL[314] WL[313] WL[312] WL[311] WL[310] WL[309] WL[308] 
+ WL[307] WL[306] WL[305] WL[304] WL[303] WL[302] WL[301] WL[300] WL[299] 
+ WL[298] WL[297] WL[296] WL[295] WL[294] WL[293] WL[292] WL[291] WL[290] 
+ WL[289] WL[288] WL[287] WL[286] WL[285] WL[284] WL[283] WL[282] WL[281] 
+ WL[280] WL[279] WL[278] WL[277] WL[276] WL[275] WL[274] WL[273] WL[272] 
+ WL[271] WL[270] WL[269] WL[268] WL[267] WL[266] WL[265] WL[264] WL[263] 
+ WL[262] WL[261] WL[260] WL[259] WL[258] WL[257] WL[256] WL[255] WL[254] 
+ WL[253] WL[252] WL[251] WL[250] WL[249] WL[248] WL[247] WL[246] WL[245] 
+ WL[244] WL[243] WL[242] WL[241] WL[240] WL[239] WL[238] WL[237] WL[236] 
+ WL[235] WL[234] WL[233] WL[232] WL[231] WL[230] WL[229] WL[228] WL[227] 
+ WL[226] WL[225] WL[224] WL[223] WL[222] WL[221] WL[220] WL[219] WL[218] 
+ WL[217] WL[216] WL[215] WL[214] WL[213] WL[212] WL[211] WL[210] WL[209] 
+ WL[208] WL[207] WL[206] WL[205] WL[204] WL[203] WL[202] WL[201] WL[200] 
+ WL[199] WL[198] WL[197] WL[196] WL[195] WL[194] WL[193] WL[192] WL[191] 
+ WL[190] WL[189] WL[188] WL[187] WL[186] WL[185] WL[184] WL[183] WL[182] 
+ WL[181] WL[180] WL[179] WL[178] WL[177] WL[176] WL[175] WL[174] WL[173] 
+ WL[172] WL[171] WL[170] WL[169] WL[168] WL[167] WL[166] WL[165] WL[164] 
+ WL[163] WL[162] WL[161] WL[160] WL[159] WL[158] WL[157] WL[156] WL[155] 
+ WL[154] WL[153] WL[152] WL[151] WL[150] WL[149] WL[148] WL[147] WL[146] 
+ WL[145] WL[144] WL[143] WL[142] WL[141] WL[140] WL[139] WL[138] WL[137] 
+ WL[136] WL[135] WL[134] WL[133] WL[132] WL[131] WL[130] WL[129] WL[128] 
+ WL[127] WL[126] WL[125] WL[124] WL[123] WL[122] WL[121] WL[120] WL[119] 
+ WL[118] WL[117] WL[116] WL[115] WL[114] WL[113] WL[112] WL[111] WL[110] 
+ WL[109] WL[108] WL[107] WL[106] WL[105] WL[104] WL[103] WL[102] WL[101] 
+ WL[100] WL[99] WL[98] WL[97] WL[96] WL[95] WL[94] WL[93] WL[92] WL[91] WL[90] 
+ WL[89] WL[88] WL[87] WL[86] WL[85] WL[84] WL[83] WL[82] WL[81] WL[80] WL[79] 
+ WL[78] WL[77] WL[76] WL[75] WL[74] WL[73] WL[72] WL[71] WL[70] WL[69] WL[68] 
+ WL[67] WL[66] WL[65] WL[64] WL[63] WL[62] WL[61] WL[60] WL[59] WL[58] WL[57] 
+ WL[56] WL[55] WL[54] WL[53] WL[52] WL[51] WL[50] WL[49] WL[48] WL[47] WL[46] 
+ WL[45] WL[44] WL[43] WL[42] WL[41] WL[40] WL[39] WL[38] WL[37] WL[36] WL[35] 
+ WL[34] WL[33] WL[32] WL[31] WL[30] WL[29] WL[28] WL[27] WL[26] WL[25] WL[24] 
+ WL[23] WL[22] WL[21] WL[20] WL[19] WL[18] WL[17] WL[16] WL[15] WL[14] WL[13] 
+ WL[12] WL[11] WL[10] WL[9] WL[8] WL[7] WL[6] WL[5] WL[4] WL[3] WL[2] WL[1] 
+ WL[0] S11000X8_TRKCOL
XCTRL AWTI BIST_BUF TIEL TIELB DCLK GW_RB WLPX WLPY WLPYB0 WLPYB1 XPD0[7] 
+ XPD0[6] XPD0[5] XPD0[4] XPD0[3] XPD0[2] XPD0[1] XPD0[0] XPD1[7] XPD1[6] 
+ XPD1[5] XPD1[4] XPD1[3] XPD1[2] XPD1[1] XPD1[0] XPD2[7] XPD2[6] XPD2[5] 
+ XPD2[4] XPD2[3] XPD2[2] XPD2[1] XPD2[0] Y10[3] Y10[2] Y10[1] Y10[0] Y32[1] 
+ Y32[0] TIELB TIELB CEB TIELB CLK TIELB TRKBL TSEL[1] TSEL[0] WEB TIELB TIELB 
+ A[11] A[10] A[9] A[8] A[7] A[6] A[5] A[4] A[3] TIELB TIELB TIELB TIELB TIELB 
+ TIELB TIELB TIELB TIELB A[2] A[1] A[0] TIELB TIELB TIELB S11000X8_CTRL888_M8
D0_0 GND A[0] NDIO 0.1066P
D0_1 GND A[1] NDIO 0.1066P
D0_2 GND A[2] NDIO 0.1066P
D0_3 GND A[3] NDIO 0.1066P
D0_4 GND A[4] NDIO 0.1066P
D0_5 GND A[5] NDIO 0.1066P
D0_6 GND A[6] NDIO 0.1066P
D0_7 GND A[7] NDIO 0.1066P
D0_8 GND A[8] NDIO 0.1066P
D0_9 GND A[9] NDIO 0.1066P
D0_10 GND A[10] NDIO 0.1066P
D0_11 GND A[11] NDIO 0.1066P
D1_0 GND D[0] NDIO 0.1066P
D10_0 GND BWEB[0] NDIO 0.1066P
D1_1 GND D[1] NDIO 0.1066P
D10_1 GND BWEB[1] NDIO 0.1066P
D1_2 GND D[2] NDIO 0.1066P
D10_2 GND BWEB[2] NDIO 0.1066P
D1_3 GND D[3] NDIO 0.1066P
D10_3 GND BWEB[3] NDIO 0.1066P
D1_4 GND D[4] NDIO 0.1066P
D10_4 GND BWEB[4] NDIO 0.1066P
D1_5 GND D[5] NDIO 0.1066P
D10_5 GND BWEB[5] NDIO 0.1066P
D1_6 GND D[6] NDIO 0.1066P
D10_6 GND BWEB[6] NDIO 0.1066P
D1_7 GND D[7] NDIO 0.1066P
D10_7 GND BWEB[7] NDIO 0.1066P
D2_CEB GND CEB NDIO 0.1066P
D3 GND CLK NDIO 0.1066P
D5 GND WEB NDIO 0.1066P
D9_0 GND TSEL[0] NDIO 0.1066P
D9_1 GND TSEL[1] NDIO 0.1066P
.ENDS

